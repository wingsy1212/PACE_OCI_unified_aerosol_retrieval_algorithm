netcdf AERDT_L2_OCI {
dimensions:
	number_of_lines_8x8 = UNLIMITED ; // e.g. 404 but varies
	number_of_pixels_8x8 = 400 ;
	number_of_lines_1x1 = UNLIMITED ; // e.g. 3232
	number_of_pixels_1x1 = 5000 ;
	Wavelength_Used_Land_1 = 3 ;
	Wavelength_Used_Land_2 = 4 ;
	Wavelength_Used_Ocean_9 = 9 ;
	Wavelength_Used_Ocean = 2 ;
    Wavelength_Used_Ocean_1 = 4 ;
	Solution_Index = 9 ;
	Quality_Flag_Num = 2 ;

// global attributes:
        :Conventions = "CF-1.6";
        :format_version = 1; 
        :instrument = "OCI";
        :platform = "";  // Suomi-NPP or NOAA-20
        :processing_level = "L2";
        :cdm_data_type = "swath";
        :creator_name = "NASA Atmosphere SIPS";
        :creator_email = "sips.support@ssec.wisc.edu";
        :creator_url = "https://sips.ssec.wisc.edu/";
        :institution = "NASA Atmosphere SIPS";
        :project = "NASA Atmosphere Discipline";
        :publisher_name = "NASA Atmosphere SIPS";
        :publisher_email = "sips.support@ssec.wisc.edu";
        :publisher_url = "https://sips.ssec.wisc.edu/";
        :keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords";
        :license = "https://science.nasa.gov/earth-science/earth-science-data/data-information-policy/";
        :stdname_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention";
        :naming_authority = "gov.nasa.gsfc.sci.atmos";
        :history = "";
        :source = "";
        :title = ""; // look this up
        :long_name = ""; // look this up
        :processing_version = "";

group: geolocation_data {
    variables:
	float longitude(number_of_lines_8x8, number_of_pixels_8x8) ;
		longitude:valid_range = -180.f, 180.f ;
		longitude:_FillValue = -999.f ;
		longitude:long_name = "Geodetic Longitude" ;
		longitude:units = "degree_east" ;
		longitude:scale_factor = 1. ;
		longitude:add_offset = 0. ;
		longitude:Parameter_Type = "OCI Input" ;
		longitude:Geolocation_Pointer = "Geolocation data not applicable" ;
		longitude:_CoordinateAxisType = "Lon" ;
        longitude:_Storage = "chunked" ;
        longitude:_ChunkSizes = 1, 400 ;
        longitude:_DeflateLevel = 5 ;
        longitude:_Shuffle = "true" ;
	float latitude(number_of_lines_8x8, number_of_pixels_8x8) ;
		latitude:valid_range = -90.f, 90.f ;
		latitude:_FillValue = -999.f ;
		latitude:long_name = "Geodetic Latitude" ;
		latitude:units = "degree_north" ;
		latitude:scale_factor = 1. ;
		latitude:add_offset = 0. ;
		latitude:Parameter_Type = "OCI Input" ;
		latitude:Geolocation_Pointer = "Geolocation data not applicable" ;
		latitude:_CoordinateAxisType = "Lat" ;
        latitude:_Storage = "chunked" ;
        latitude:_ChunkSizes = 1, 400 ;
        latitude:_DeflateLevel = 5 ;
        latitude:_Shuffle = "true" ;
	short solar_zenith_angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		solar_zenith_angle:valid_range = 0s, 18000s ;
		solar_zenith_angle:_FillValue = -9999s ;
		solar_zenith_angle:long_name = "Solar Zenith Angle, Cell to Sun" ;
		solar_zenith_angle:units = "degree" ;
		solar_zenith_angle:scale_factor = 0.01 ;
		solar_zenith_angle:add_offset = 0. ;
		solar_zenith_angle:Parameter_Type = "OCI Input" ;
		solar_zenith_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		solar_zenith_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        solar_zenith_angle:_Storage = "chunked" ;
        solar_zenith_angle:_ChunkSizes = 1, 400 ;
        solar_zenith_angle:_DeflateLevel = 5 ;
        solar_zenith_angle:_Shuffle = "true" ;
	short solar_azimuth_angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		solar_azimuth_angle:valid_range = -18000s, 18000s ;
		solar_azimuth_angle:_FillValue = -9999s ;
		solar_azimuth_angle:long_name = "Solar Azimuth Angle, Cell to Sun" ;
		solar_azimuth_angle:units = "degree" ;
		solar_azimuth_angle:scale_factor = 0.01 ;
		solar_azimuth_angle:add_offset = 0. ;
		solar_azimuth_angle:Parameter_Type = "OCI Input" ;
		solar_azimuth_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		solar_azimuth_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        solar_azimuth_angle:_Storage = "chunked" ;
        solar_azimuth_angle:_ChunkSizes = 1, 400 ;
        solar_azimuth_angle:_DeflateLevel = 5 ;
        solar_azimuth_angle:_Shuffle = "true" ;
	short sensor_zenith_angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		sensor_zenith_angle:valid_range = 0s, 18000s ;
		sensor_zenith_angle:_FillValue = -9999s ;
		sensor_zenith_angle:long_name = "Sensor Zenith Angle, Cell to Sensor" ;
		sensor_zenith_angle:units = "degree" ;
		sensor_zenith_angle:scale_factor = 0.01 ;
		sensor_zenith_angle:add_offset = 0. ;
		sensor_zenith_angle:Parameter_Type = "OCI Input" ;
		sensor_zenith_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		sensor_zenith_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        sensor_zenith_angle:_Storage = "chunked" ;
        sensor_zenith_angle:_ChunkSizes = 1, 400 ;
        sensor_zenith_angle:_DeflateLevel = 5 ;
        sensor_zenith_angle:_Shuffle = "true" ;
	short sensor_azimuth_angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		sensor_azimuth_angle:valid_range = -18000s, 18000s ;
		sensor_azimuth_angle:_FillValue = -9999s ;
		sensor_azimuth_angle:long_name = "Sensor Azimuth Angle, Cell to Sensor" ;
		sensor_azimuth_angle:units = "degree" ;
		sensor_azimuth_angle:scale_factor = 0.01 ;
		sensor_azimuth_angle:add_offset = 0. ;
		sensor_azimuth_angle:Parameter_Type = "OCI Input" ;
		sensor_azimuth_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		sensor_azimuth_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        sensor_azimuth_angle:_Storage = "chunked" ;
        sensor_azimuth_angle:_ChunkSizes = 1, 400 ;
        sensor_azimuth_angle:_DeflateLevel = 5 ;
        sensor_azimuth_angle:_Shuffle = "true" ; 
    data:
    } // group geolocation_data
group: geophysical_data {
    variables:
	short Effective_Optical_Depth_Average_Ocean_UV(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean_9) ;
		Effective_Optical_Depth_Average_Ocean_UV:valid_range = -50s, 5000s ;
		Effective_Optical_Depth_Average_Ocean_UV:_FillValue = -9999s ;
		Effective_Optical_Depth_Average_Ocean_UV:long_name = "Retrieved AOT for 0.354,0.388 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Effective_Optical_Depth_Average_Ocean_UV:units = "None" ;
		Effective_Optical_Depth_Average_Ocean_UV:scale_factor = 0.001 ;
		Effective_Optical_Depth_Average_Ocean_UV:add_offset = 0. ;
		Effective_Optical_Depth_Average_Ocean_UV:Parameter_Type = "Output" ;
		Effective_Optical_Depth_Average_Ocean_UV:Geolocation_Pointer = "Internal geolocation arrays" ;
		Effective_Optical_Depth_Average_Ocean_UV:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Effective_Optical_Depth_Average_Ocean_UV:_Storage = "chunked" ;
        Effective_Optical_Depth_Average_Ocean_UV:_ChunkSizes = 1, 400, 4 ;
        Effective_Optical_Depth_Average_Ocean_UV:_DeflateLevel = 5 ;
        Effective_Optical_Depth_Average_Ocean_UV:_Shuffle = "true" ;
	
       short Single_Scattering_Albedo_Average_Ocean_UV(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		Single_Scattering_Albedo_Average_Ocean_UV:valid_range = 700s, 1000s ;
		Single_Scattering_Albedo_Average_Ocean_UV:_FillValue = -9999s ;
		Single_Scattering_Albedo_Average_Ocean_UV:long_name = "Single scattering Albedo  0.354 and 0.388 microns" ;
		Single_Scattering_Albedo_Average_Ocean_UV:units = "None" ;
		Single_Scattering_Albedo_Average_Ocean_UV:scale_factor = 0.001 ;
		Single_Scattering_Albedo_Average_Ocean_UV:add_offset = 0. ;
		Single_Scattering_Albedo_Average_Ocean_UV:Parameter_Type = "Output" ;
		Single_Scattering_Albedo_Average_Ocean_UV:Geolocation_Pointer = "Internal geolocation arrays" ;
		Single_Scattering_Albedo_Average_Ocean_UV:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        
   short Optical_Depth_Ratio_Small_Ocean_used(number_of_lines_8x8, number_of_pixels_8x8) ;
		Optical_Depth_Ratio_Small_Ocean_used:valid_range = 0s, 1000s ;
		Optical_Depth_Ratio_Small_Ocean_used:_FillValue = -9999s ;
		Optical_Depth_Ratio_Small_Ocean_used:long_name = "Fraction of AOT (at 0.55 micron) contributed by fine mode used for UV retrieval" ;
		Optical_Depth_Ratio_Small_Ocean_used:units = "None" ;
		Optical_Depth_Ratio_Small_Ocean_used:scale_factor = 0.001 ;
		Optical_Depth_Ratio_Small_Ocean_used:add_offset = 0. ;
		Optical_Depth_Ratio_Small_Ocean_used:Parameter_Type = "Output" ;
		Optical_Depth_Ratio_Small_Ocean_used:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Ratio_Small_Ocean_used:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Optical_Depth_Ratio_Small_Ocean_used:_Storage = "chunked" ;
        Optical_Depth_Ratio_Small_Ocean_used:_ChunkSizes = 1, 400 ;
        Optical_Depth_Ratio_Small_Ocean_used:_DeflateLevel = 5 ;
        Optical_Depth_Ratio_Small_Ocean_used:_Shuffle = "true" ;
    short Fine_MODE_used(number_of_lines_8x8, number_of_pixels_8x8) ;
		Fine_MODE_used:valid_range = 1s, 4s ;
		Fine_MODE_used:_FillValue = -9999s ;
		Fine_MODE_used:long_name = "Fine MODE used for  UV retrieval " ;
		Fine_MODE_used:units = "Meters/sec" ;
		Fine_MODE_used:scale_factor = 1 ;
		Fine_MODE_used:add_offset = 0. ;
		Fine_MODE_used:Parameter_Type = "Output" ;
		Fine_MODE_used:Geolocation_Pointer = "Internal geolocation arrays" ;
		Fine_MODE_used:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Fine_MODE_used:_Storage = "chunked" ;
        Fine_MODE_used:_ChunkSizes = 1, 400 ;
        Fine_MODE_used:_DeflateLevel = 5 ;
        Fine_MODE_used:_Shuffle = "true" ;
    short Coarse_MODE_used(number_of_lines_8x8, number_of_pixels_8x8) ;
		Coarse_MODE_used:valid_range = 1s, 6s ;
		Coarse_MODE_used:_FillValue = -9999s ;
		Coarse_MODE_used:long_name = "Coarse MODE used for UV retrieval ";
		Coarse_MODE_used:units = "None" ;
		Coarse_MODE_used:scale_factor = 1 ;
		Coarse_MODE_used:add_offset = 0. ;
		Coarse_MODE_used:Parameter_Type = "Output" ;
		Coarse_MODE_used:Geolocation_Pointer = "Internal geolocation arrays" ;
		Coarse_MODE_used:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Coarse_MODE_used:_Storage = "chunked" ;
        Coarse_MODE_used:_ChunkSizes = 1, 400 ;
        Coarse_MODE_used:_DeflateLevel = 5 ;
        Coarse_MODE_used:_Shuffle = "true" ;
      short Index_Albedo(number_of_lines_8x8, number_of_pixels_8x8) ;
		Index_Albedo:valid_range = 1s, 4s ;
		Index_Albedo:_FillValue = -9999s ;
		Index_Albedo:long_name = "Index for Single scattering Albedo1=nabsor,2=dust,3=C1,4=C2";
		Index_Albedo:units = "None" ;
		Index_Albedo:scale_factor = 1 ;
		Index_Albedo:add_offset = 0. ;
		Index_Albedo:Parameter_Type = "Output" ;
		Index_Albedo:Geolocation_Pointer = "Internal geolocation arrays" ;
		Index_Albedo:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Index_Albedo:_Storage = "chunked" ;
        Index_Albedo:_ChunkSizes = 1, 400 ;
        Index_Albedo:_DeflateLevel = 5 ;
        Index_Albedo:_Shuffle = "true" ;
     short Height(number_of_lines_8x8, number_of_pixels_8x8) ;
		Height:valid_range = 1s, 10s ;
		Height:_FillValue = -9999s ;
		Height:long_name = "Height 1.5KM  3KM, 6KM, 10KM)";
		Height:units = "KM" ;
		Height:scale_factor = 1 ;
		Height:add_offset = 0. ;
		Height:Parameter_Type = "Output" ;
		Height:Geolocation_Pointer = "Internal geolocation arrays" ;
		Height:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Height:_Storage = "chunked" ;
        Height:_ChunkSizes = 1, 400 ;
        Height:_DeflateLevel = 5 ;
        Height:_Shuffle = "true" ;
      short Fitting_Error_Height(number_of_lines_8x8, number_of_pixels_8x8) ;
		Fitting_Error_Height:valid_range = 0s, 10000s ;
		Fitting_Error_Height:_FillValue = -9999s ;
		Fitting_Error_Height:long_name = "Fitting_Error_Height" ;
		Fitting_Error_Height:units = "None" ;
		Fitting_Error_Height:scale_factor = 0.001 ;
		Fitting_Error_Height:add_offset = 0. ;
		Fitting_Error_Height:Parameter_Type = "Output" ;
		Fitting_Error_Height:Geolocation_Pointer = "Internal geolocation arrays" ;
		Fitting_Error_Height:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Fitting_Error_Height:_Storage = "chunked" ;
        Fitting_Error_Height:_ChunkSizes = 1, 400 ;
        Fitting_Error_Height:_DeflateLevel = 5 ;
        Fitting_Error_Height:_Shuffle = "true" ;
        short Mean_Reflectance_UV_ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean_9) ;
		Mean_Reflectance_UV_ocean:valid_range = 0s, 10000s ;
		Mean_Reflectance_UV_ocean:_FillValue = -9999s ;
		Mean_Reflectance_UV_ocean:long_name = "Mean reflectance of pixels used for Ocean 0.354,0.388 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Mean_Reflectance_UV_ocean:units = "None" ;
		Mean_Reflectance_UV_ocean:scale_factor = 0.0001 ;
		Mean_Reflectance_UV_ocean:add_offset = 0. ;
		Mean_Reflectance_UV_ocean:Parameter_Type = "Output" ;
		Mean_Reflectance_UV_ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mean_Reflectance_UV_ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		
    data:
    } // group geophysical_data
}

