netcdf AERDT_L2_OCI {
dimensions:
	number_of_lines_7x7 = UNLIMITED ; // e.g. 404 but varies
	number_of_pixels_7x7 = 181 ;
	Wavelength_Used_all = 9 ; 
	Wavelength_Used_DTDB = 7 ; 
	Wavelength_Used_UV = 3 ; 
	Wavelength_Used_UV1 = 2 ;
	Wavelength_ACA_UNCER = 2 ;
	Wavelength_Used = 5 ;
	Height_Levels = 5;
	
// global attributes:
        :Conventions = "CF-1.6";
        :format_version = 1; 
        :instrument = "OCI";
        :platform = "";  // Suomi-NPP or NOAA-20
        :processing_level = "L2";
        :cdm_data_type = "swath";
        :creator_name = "NASA Atmosphere SIPS";
        :creator_email = "sips.support@ssec.wisc.edu";
        :creator_url = "https://sips.ssec.wisc.edu/";
        :institution = "NASA Atmosphere SIPS";
        :project = "NASA Atmosphere Discipline";
        :publisher_name = "NASA Atmosphere SIPS";
        :publisher_email = "sips.support@ssec.wisc.edu";
        :publisher_url = "https://sips.ssec.wisc.edu/";
        :keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords";
        :license = "https://science.nasa.gov/earth-science/earth-science-data/data-information-policy/";
        :stdname_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention";
        :naming_authority = "gov.nasa.gsfc.sci.atmos";
        :history = "";
        :source = "";
        :title = ""; // look this up
        :long_name = ""; // look this up
        :processing_version = "";

group: geolocation_data {
    variables:
	
	float longitude(number_of_lines_7x7, number_of_pixels_7x7) ;
		longitude:valid_range = -180.f, 180.f ;
		longitude:_FillValue = -999.f ;
		longitude:long_name = "Geodetic Longitude" ;
		longitude:units = "degree_east" ;
		longitude:scale_factor = 1. ;
		longitude:add_offset = 0. ;
		longitude:Parameter_Type = "OCI Input" ;
		longitude:Geolocation_Pointer = "Geolocation data not applicable" ;
		longitude:_CoordinateAxisType = "Lon" ;
		longitude:_ChunkSizes = 32, 32 ;
		longitude:_DeflateLevel = 4 ;
         
	float latitude(number_of_lines_7x7, number_of_pixels_7x7) ;
		latitude:valid_range = -90.f, 90.f ;
		latitude:_FillValue = -999.f ;
		latitude:long_name = "Geodetic Latitude" ;
		latitude:units = "degree_north" ;
		latitude:scale_factor = 1. ;
		latitude:add_offset = 0. ;
		latitude:Parameter_Type = "OCI Input" ;
		latitude:Geolocation_Pointer = "Geolocation data not applicable" ;
		latitude:_CoordinateAxisType = "Lat" ;
		latitude:_ChunkSizes = 32, 32 ;
 		latitude:_DeflateLevel = 4 ;
         
	short solar_zenith_angle(number_of_lines_7x7, number_of_pixels_7x7) ;
		solar_zenith_angle:valid_range = 0s, 18000s ;
		solar_zenith_angle:_FillValue = -9999s ;
		solar_zenith_angle:long_name = "Solar Zenith Angle, Cell to Sun" ;
		solar_zenith_angle:units = "degree" ;
		solar_zenith_angle:scale_factor = 0.01 ;
		solar_zenith_angle:add_offset = 0. ;
		solar_zenith_angle:Parameter_Type = "OCI Input" ;
		solar_zenith_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		solar_zenith_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		solar_azimuth_angle:_ChunkSizes = 32, 32 ;
		solar_zenith_angle:_DeflateLevel = 4 ;
         
	short solar_azimuth_angle(number_of_lines_7x7, number_of_pixels_7x7) ;
		solar_azimuth_angle:valid_range = -18000s, 18000s ;
		solar_azimuth_angle:_FillValue = -9999s ;
		solar_azimuth_angle:long_name = "Solar Azimuth Angle, Cell to Sun" ;
		solar_azimuth_angle:units = "degree" ;
		solar_azimuth_angle:scale_factor = 0.01 ;
		solar_azimuth_angle:add_offset = 0. ;
		solar_azimuth_angle:Parameter_Type = "OCI Input" ;
		solar_azimuth_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		solar_azimuth_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		solar_azimuth_angle:_ChunkSizes = 32, 32 ;
		solar_azimuth_angle:_DeflateLevel = 4 ;
         
	short sensor_zenith_angle(number_of_lines_7x7, number_of_pixels_7x7) ;
		sensor_zenith_angle:valid_range = 0s, 18000s ;
		sensor_zenith_angle:_FillValue = -9999s ;
		sensor_zenith_angle:long_name = "Sensor Zenith Angle, Cell to Sensor" ;
		sensor_zenith_angle:units = "degree" ;
		sensor_zenith_angle:scale_factor = 0.01 ;
		sensor_zenith_angle:add_offset = 0. ;
		sensor_zenith_angle:Parameter_Type = "OCI Input" ;
		sensor_zenith_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		sensor_zenith_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		sensor_zenith_angle:_ChunkSizes = 32, 32 ;
		sensor_zenith_angle:_DeflateLevel = 4 ;
        
	short sensor_azimuth_angle(number_of_lines_7x7, number_of_pixels_7x7) ;
		sensor_azimuth_angle:valid_range = -18000s, 18000s ;
		sensor_azimuth_angle:_FillValue = -9999s ;
		sensor_azimuth_angle:long_name = "Sensor Azimuth Angle, Cell to Sensor" ;
		sensor_azimuth_angle:units = "degree" ;
		sensor_azimuth_angle:scale_factor = 0.01 ;
		sensor_azimuth_angle:add_offset = 0. ;
		sensor_azimuth_angle:Parameter_Type = "OCI Input" ;
		sensor_azimuth_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		sensor_azimuth_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		sensor_azimuth_angle:_ChunkSizes = 32, 32 ;
		sensor_azimuth_angle:_DeflateLevel = 4 ;
        
    data:
    } // group geolocation_data

group: geophysical_data {
    variables:
   short Land_Sea_Flag(number_of_lines_7x7, number_of_pixels_7x7) ;
		Land_Sea_Flag:valid_range = 0s, 1s ;
		Land_Sea_Flag:_FillValue = -9999s ;
		Land_Sea_Flag:long_name = "Land_Sea_Flag( 0 = Ocean, 1 = Land )" ;
		Land_Sea_Flag:units = "None" ;
		Land_Sea_Flag:scale_factor = 1. ;
		Land_Sea_Flag:add_offset = 0. ;
		Land_Sea_Flag:Parameter_Type = "Output" ;
		Land_Sea_Flag:Geolocation_Pointer = "Internal geolocation arrays" ;
		Land_Sea_Flag:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		Land_Sea_Flag:_ChunkSizes = 32, 32 ;
		Land_Sea_Flag:_DeflateLevel = 4 ;
                 
   short Aerosol_Optical_Depth(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_Used_all) ;
		Aerosol_Optical_Depth:valid_range = -50s, 5000s ;
		Aerosol_Optical_Depth:_FillValue = -9999s ;
		Aerosol_Optical_Depth:long_name = "Retrieved AOT at 0.354,0.388 0.48, 0.55, 0.67, 0.87 1.24, 1.64, 2.2"  ;
		Aerosol_Optical_Depth:units = "None" ;
		Aerosol_Optical_Depth:scale_factor = 0.001 ;
		Aerosol_Optical_Depth:add_offset = 0. ;
		Aerosol_Optical_Depth:Parameter_Type = "Output" ;
		Aerosol_Optical_Depth:Geolocation_Pointer = "Internal geolocation arrays" ;
		Aerosol_Optical_Depth:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		Aerosol_Optical_Depth:_ChunkSizes = 32, 32, 9 ;
		Aerosol_Optical_Depth:_DeflateLevel = 4 ;
         
   short Optical_Depth_Ratio_Small_Ocean_used(number_of_lines_7x7, number_of_pixels_7x7) ;
		Optical_Depth_Ratio_Small_Ocean_used:valid_range = 0s, 1000s ;
		Optical_Depth_Ratio_Small_Ocean_used:_FillValue = -9999s ;
		Optical_Depth_Ratio_Small_Ocean_used:long_name = "Fraction of AOT (at 0.55 micron) contributed by fine mode used for UV retrieval" ;
		Optical_Depth_Ratio_Small_Ocean_used:units = "None" ;
		Optical_Depth_Ratio_Small_Ocean_used:scale_factor = 0.001 ;
		Optical_Depth_Ratio_Small_Ocean_used:add_offset = 0. ;
		Optical_Depth_Ratio_Small_Ocean_used:Parameter_Type = "Output" ;
		Optical_Depth_Ratio_Small_Ocean_used:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Ratio_Small_Ocean_used:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		Optical_Depth_Ratio_Small_Ocean_used:_ChunkSizes = 32, 32 ;
		Optical_Depth_Ratio_Small_Ocean_used:_DeflateLevel = 4 ;
             
   short Mean_Gas_Corrected_Reflectance(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_Used_DTDB) ;
		Mean_Gas_Corrected_Reflectance:valid_range = 0s, 10000s ;
		Mean_Gas_Corrected_Reflectance:_FillValue = -9999s ;
		Mean_Gas_Corrected_Reflectance:long_name = "Mean reflectance Gas corrected of pixels at  0.48, 0.55, 0.67, 0.87 1.24, 1.64, 2.2" ;
		Mean_Gas_Corrected_Reflectance:units = "None" ;
		Mean_Gas_Corrected_Reflectance:scale_factor = 0.0001 ;
		Mean_Gas_Corrected_Reflectance:add_offset = 0. ;
		Mean_Gas_Corrected_Reflectance:Parameter_Type = "Output" ;
		Mean_Gas_Corrected_Reflectance:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mean_Gas_Corrected_Reflectance:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		Mean_Gas_Corrected_Reflectance:_ChunkSizes = 32, 32, 7 ;
		Mean_Gas_Corrected_Reflectance:_DeflateLevel = 4 ;
		
  short Mean_Reflectance(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_Used_UV1);
		Mean_Reflectance:valid_range = 0s, 10000s ;
		Mean_Reflectance:_FillValue = -9999s ;
		Mean_Reflectance:long_name = "Mean reflectance (not corrected for GAS ) pixels at 0.354 0.388" ;
		Mean_Reflectance:units = "None" ;
		Mean_Reflectance:scale_factor = 0.0001 ;
		Mean_Reflectance:add_offset = 0. ;
		Mean_Reflectance:Parameter_Type = "Output" ;
		Mean_Reflectance:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mean_Reflectance:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		Mean_Reflectance:_ChunkSizes = 32, 32, 2 ;
		Mean_Reflectance:_DeflateLevel = 4 ;
       
    short  DT_AerosolSingleScattAlbedo(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_Used_UV) ;
		DT_AerosolSingleScattAlbedo:valid_range = 700s, 1000s ;
		DT_AerosolSingleScattAlbedo:_FillValue = -9999s ;
		DT_AerosolSingleScattAlbedo:long_name = "Single scattering Albedo from Dark Target ocean 0.354 and 0.388 and 0.50, microns" ;
		DT_AerosolSingleScattAlbedo:units = "None" ;
		DT_AerosolSingleScattAlbedo:scale_factor = 0.001 ;
		DT_AerosolSingleScattAlbedo:add_offset = 0. ;
		DT_AerosolSingleScattAlbedo:Parameter_Type = "Output" ;
		DT_AerosolSingleScattAlbedo:Geolocation_Pointer = "Internal geolocation arrays" ;
		DT_AerosolSingleScattAlbedo:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;	
		DT_AerosolSingleScattAlbedo:_ChunkSizes = 32, 32, 3 ;
		DT_AerosolSingleScattAlbedo:_DeflateLevel = 4 ;
		
    short DT_AerosolLayerHeight(number_of_lines_7x7, number_of_pixels_7x7) ;
		DT_AerosolLayerHeight:valid_range = 1s, 10s ;
		DT_AerosolLayerHeight:_FillValue = -9999s ;
		DT_AerosolLayerHeight:long_name = "Height 1.5KM  3KM, 6KM, 10KM)";
		DT_AerosolLayerHeight:units = "KM" ;
		DT_AerosolLayerHeight:scale_factor = 1 ;
		DT_AerosolLayerHeight:add_offset = 0. ;
		DT_AerosolLayerHeight:Parameter_Type = "Output" ;
		DT_AerosolLayerHeight:Geolocation_Pointer = "Internal geolocation arrays" ;
		DT_AerosolLayerHeight:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		DT_AerosolLayerHeight:_ChunkSizes = 32, 32 ;
		DT_AerosolLayerHeight:_DeflateLevel = 4 ;
        
    short Aerosol_Cld_Fraction_Land_Ocean(number_of_lines_7x7, number_of_pixels_7x7) ;
		Aerosol_Cld_Fraction_Land_Ocean:valid_range = 0S, 1000S ;
		Aerosol_Cld_Fraction_Land_Ocean:_FillValue = -9999s ;
		Aerosol_Cld_Fraction_Land_Ocean:long_name = "Aerosol Cloud Fraction in each box" ;
		Aerosol_Cld_Fraction_Land_Ocean:units = "None" ;
		Aerosol_Cld_Fraction_Land_Ocean:scale_factor = 0.001 ;
		Aerosol_Cld_Fraction_Land_Ocean:add_offset = 0. ;
		Aerosol_Cld_Fraction_Land_Ocean:Parameter_Type = "Output" ;
		Aerosol_Cld_Fraction_Land_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Aerosol_Cld_Fraction_Land_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		Aerosol_Cld_Fraction_Land_Ocean:_ChunkSizes = 32, 32 ;
		Aerosol_Cld_Fraction_Land_Ocean:_DeflateLevel = 4 ;

	short NUV_AerosolIndex(number_of_lines_7x7, number_of_pixels_7x7) ;
		NUV_AerosolIndex:valid_range =  -5000s, 10000s ; 
		NUV_AerosolIndex:_FillValue = -9999s ;
		NUV_AerosolIndex:long_name = "NUV Retrieved Aerosol Index (0.354,0.388) Pair"  ;
		NUV_AerosolIndex:units = "None" ;
		NUV_AerosolIndex:scale_factor = 0.001 ;
		NUV_AerosolIndex:add_offset = 0. ;
		NUV_AerosolIndex:Parameter_Type = "Output" ;
		NUV_AerosolIndex:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_AerosolIndex:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;  
		NUV_AerosolIndex:_ChunkSizes = 32, 32 ;
		NUV_AerosolIndex:_DeflateLevel = 4 ;
	      
	short NUV_AerosolLayerHeight(number_of_lines_7x7, number_of_pixels_7x7) ;
		NUV_AerosolLayerHeight:valid_range = 0s, 10000s ;
		NUV_AerosolLayerHeight:_FillValue = -9999s ;
		NUV_AerosolLayerHeight:long_name = "NUV Retrieved Aerosol Layer Height";
		NUV_AerosolLayerHeight:units = "km" ;
		NUV_AerosolLayerHeight:scale_factor = 0.001 ;
		NUV_AerosolLayerHeight:add_offset = 0. ;
		NUV_AerosolLayerHeight:Parameter_Type = "Output" ;
		NUV_AerosolLayerHeight:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_AerosolLayerHeight:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;  
		NUV_AerosolLayerHeight:_ChunkSizes = 32, 32 ;
		NUV_AerosolLayerHeight:_DeflateLevel = 4 ;
		
	short NUV_AerosolSingleScattAlbedo(number_of_lines_7x7, number_of_pixels_7x7,Wavelength_Used) ;
		NUV_AerosolSingleScattAlbedo:valid_range = 700s, 1000s ;
		NUV_AerosolSingleScattAlbedo:_FillValue = -9999s ;
		NUV_AerosolSingleScattAlbedo:long_name = "NUV Retrieved Aerosol Single Scattering Albedo at 0.354, 0.388, 0.480, 0.550, 0.670" ;
		NUV_AerosolSingleScattAlbedo:units = "None" ;
		NUV_AerosolSingleScattAlbedo:scale_factor = 0.001 ;
		NUV_AerosolSingleScattAlbedo:add_offset = 0. ;
		NUV_AerosolSingleScattAlbedo:Parameter_Type = "Output" ;
		NUV_AerosolSingleScattAlbedo:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_AerosolSingleScattAlbedo:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;	
		NUV_AerosolSingleScattAlbedo:_ChunkSizes = 32, 32, 5 ;
		NUV_AerosolSingleScattAlbedo:_DeflateLevel = 4 ;
        
	short NUV_RadiativeCloudFraction(number_of_lines_7x7, number_of_pixels_7x7) ;
		NUV_RadiativeCloudFraction:valid_range = 0s, 1000s ;
		NUV_RadiativeCloudFraction:_FillValue = -9999s ;
		NUV_RadiativeCloudFraction:long_name = "NUV derived Radiative Equivalent Cloud Fraction at 0.388"  ;
		NUV_RadiativeCloudFraction:units = "None" ;
		NUV_RadiativeCloudFraction:scale_factor = 0.001;
		NUV_RadiativeCloudFraction:add_offset = 0. ;
		NUV_RadiativeCloudFraction:Parameter_Type = "Output" ;
		NUV_RadiativeCloudFraction:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_RadiativeCloudFraction:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_RadiativeCloudFraction:_ChunkSizes = 32, 32 ;
		NUV_RadiativeCloudFraction:_DeflateLevel = 4 ;
         
	short NUV_Residue(number_of_lines_7x7, number_of_pixels_7x7) ;
		NUV_Residue:valid_range = -5000s, 10000s ;
		NUV_Residue:_FillValue = -9999s ;
		NUV_Residue:long_name = "NUV Retrieved LER based AI (0.354,0.388) Pair"  ;
		NUV_Residue:units = "None" ;
		NUV_Residue:scale_factor = 0.001 ;
		NUV_Residue:add_offset = 0. ;
		NUV_Residue:Parameter_Type = "Output" ;
		NUV_Residue:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_Residue:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_Residue:_ChunkSizes = 32, 32 ;
		NUV_Residue:_DeflateLevel = 4 ;

	short NUV_Reflectivity(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_Used_UV1) ;
		NUV_Reflectivity:valid_range = 0s, 1000s ;
		NUV_Reflectivity:_FillValue = -9999s ;
		NUV_Reflectivity:long_name = "NUV Retrieved Aerosol Optical Depth Over Cloud at 0.354, 0.388"  ;
		NUV_Reflectivity:units = "None" ;
		NUV_Reflectivity:scale_factor = 0.001 ;
		NUV_Reflectivity:add_offset = 0.0 ;
		NUV_Reflectivity:Parameter_Type = "Output" ;
		NUV_Reflectivity:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_Reflectivity:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_Reflectivity:_ChunkSizes = 32, 32, 2 ;
		NUV_Reflectivity:_DeflateLevel = 4 ;

	short NUV_CloudOpticalDepth(number_of_lines_7x7, number_of_pixels_7x7) ;
		NUV_CloudOpticalDepth:valid_range = 0s, 5000s ;
		NUV_CloudOpticalDepth:_FillValue = -9999s ;
		NUV_CloudOpticalDepth:long_name = "NUV Retrieved Cloud Optical Depth at 0.388"  ;
		NUV_CloudOpticalDepth:units = "None" ;
		NUV_CloudOpticalDepth:scale_factor = 0.001 ;
		NUV_CloudOpticalDepth:add_offset = 0. ;
		NUV_CloudOpticalDepth:Parameter_Type = "Output" ;
		NUV_CloudOpticalDepth:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_CloudOpticalDepth:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_CloudOpticalDepth:_ChunkSizes = 32, 32 ;
		NUV_CloudOpticalDepth:_DeflateLevel = 4 ;
         
	short NUV_AerosolOpticalDepthOverCloud(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_Used_UV) ;
		NUV_AerosolOpticalDepthOverCloud:valid_range = 0s, 5000s ;
		NUV_AerosolOpticalDepthOverCloud:_FillValue = -9999s ;
		NUV_AerosolOpticalDepthOverCloud:long_name = "NUV Retrieved Aerosol Optical Depth Over Cloud at 0.354, 0.388, 0.550"  ;
		NUV_AerosolOpticalDepthOverCloud:units = "None" ;
		NUV_AerosolOpticalDepthOverCloud:scale_factor = 0.001 ;
		NUV_AerosolOpticalDepthOverCloud:add_offset = 0.0 ;
		NUV_AerosolOpticalDepthOverCloud:Parameter_Type = "Output" ;
		NUV_AerosolOpticalDepthOverCloud:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_AerosolOpticalDepthOverCloud:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_AerosolOpticalDepthOverCloud:_ChunkSizes = 32, 32, 3 ;
		NUV_AerosolOpticalDepthOverCloud:_DeflateLevel = 4 ;
         
	short NUV_AerosolCorrCloudOpticalDepth(number_of_lines_7x7, number_of_pixels_7x7) ;
		NUV_AerosolCorrCloudOpticalDepth:valid_range = 0s, 500s ;
		NUV_AerosolCorrCloudOpticalDepth:_FillValue = -9999s ;
		NUV_AerosolCorrCloudOpticalDepth:long_name = "NUV Retrieved Aerosol Corrected Cloud Optical Depth at 0.388"  ;
		NUV_AerosolCorrCloudOpticalDepth:units = "None" ;
		NUV_AerosolCorrCloudOpticalDepth:scale_factor = 0.1 ;
		NUV_AerosolCorrCloudOpticalDepth:add_offset = 0. ;
		NUV_AerosolCorrCloudOpticalDepth:Parameter_Type = "Output" ;
		NUV_AerosolCorrCloudOpticalDepth:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_AerosolCorrCloudOpticalDepth:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_AerosolCorrCloudOpticalDepth:_ChunkSizes = 32, 32 ;
		NUV_AerosolCorrCloudOpticalDepth:_DeflateLevel = 4 ;

	short NUV_AerosolOpticalDepthOverCloudVsHeight(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_Used_UV, Height_Levels) ;
		NUV_AerosolOpticalDepthOverCloud:valid_range = 0s, 5000s ;
		NUV_AerosolOpticalDepthOverCloud:_FillValue = -9999s ;
		NUV_AerosolOpticalDepthOverCloud:long_name = "NUV Retrieved Aerosol Optical Depth Over Cloud for 0.354, 0.388, 0.550 at 5 levels"  ;
		NUV_AerosolOpticalDepthOverCloud:units = "None" ;
		NUV_AerosolOpticalDepthOverCloud:scale_factor = 0.001 ;
		NUV_AerosolOpticalDepthOverCloud:add_offset = 0.0 ;
		NUV_AerosolOpticalDepthOverCloud:Parameter_Type = "Output" ;
		NUV_AerosolOpticalDepthOverCloud:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_AerosolOpticalDepthOverCloud:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_AerosolOpticalDepthOverCloud:_ChunkSizes = 32, 32, 3, 5 ;
		NUV_AerosolOpticalDepthOverCloud:_DeflateLevel = 4 ;
         
	short NUV_AerosolCorrCloudOpticalDepthVsHeight(number_of_lines_7x7, number_of_pixels_7x7, Height_Levels) ;
		NUV_AerosolCorrCloudOpticalDepth:valid_range = 0s, 500s ;
		NUV_AerosolCorrCloudOpticalDepth:_FillValue = -9999s ;
		NUV_AerosolCorrCloudOpticalDepth:long_name = "NUV Retrieved Aerosol Corrected Cloud Optical Depth for 0.388 micron at 5 levels"  ;
		NUV_AerosolCorrCloudOpticalDepth:units = "None" ;
		NUV_AerosolCorrCloudOpticalDepth:scale_factor = 0.1 ;
		NUV_AerosolCorrCloudOpticalDepth:add_offset = 0. ;
		NUV_AerosolCorrCloudOpticalDepth:Parameter_Type = "Output" ;
		NUV_AerosolCorrCloudOpticalDepth:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_AerosolCorrCloudOpticalDepth:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_AerosolCorrCloudOpticalDepth:_ChunkSizes = 32, 32, 5 ;
		NUV_AerosolCorrCloudOpticalDepth:_DeflateLevel = 4 ;

	short NUV_FinalAlgorithmFlagsACA(number_of_lines_7x7, number_of_pixels_7x7) ;
		NUV_FinalAlgorithmFlagsACA:valid_range = 0s, 3000s ;
		NUV_FinalAlgorithmFlagsACA:_FillValue = -9999s ;
		NUV_FinalAlgorithmFlagsACA:long_name = "NUV Final Algorithm Flags for Above-cloud retrievals"  ;
		NUV_FinalAlgorithmFlagsACA:units = "None" ;
		NUV_FinalAlgorithmFlagsACA:scale_factor = 0.001 ;
		NUV_FinalAlgorithmFlagsACA:add_offset = 0. ;
		NUV_FinalAlgorithmFlagsACA:Parameter_Type = "Output" ;
		NUV_FinalAlgorithmFlagsACA:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_FinalAlgorithmFlagsACA:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_FinalAlgorithmFlagsACA:_ChunkSizes = 32, 32 ;
		NUV_FinalAlgorithmFlagsACA:_DeflateLevel = 4 ;

	short NUV_UncertaintyACAODToSSA(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_ACA_UNCER) ;
		NUV_UncertaintyACAODToSSA:valid_range = -1000s, 1000s ;
		NUV_UncertaintyACAODToSSA:_FillValue = -9999s ;
		NUV_UncertaintyACAODToSSA:long_name = "NUV derived percent uncertainity in COD due to change in SSA." ;
		NUV_UncertaintyACAODToSSA:units = "None" ;
		NUV_UncertaintyACAODToSSA:scale_factor = 0.1 ;
		NUV_UncertaintyACAODToSSA:add_offset = 0. ;
		NUV_UncertaintyACAODToSSA:Parameter_Type = "Output" ;
		NUV_UncertaintyACAODToSSA:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_UncertaintyACAODToSSA:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_UncertaintyACAODToSSA:_ChunkSizes = 32, 32, 2 ;
		NUV_UncertaintyACAODToSSA:_DeflateLevel = 4 ;
		
	short NUV_UncertaintyCODToSSA(number_of_lines_7x7, number_of_pixels_7x7, Wavelength_ACA_UNCER) ;
		NUV_UncertaintyCODToSSA:valid_range = -1000s, 1000s ;
		NUV_UncertaintyCODToSSA:_FillValue = -9999s ;
		NUV_UncertaintyCODToSSA:long_name = "NUV derived percent uncertainity in Aerosol-corrected COD due to plus/minus 0.03 change in SSA."  ;
		NUV_UncertaintyCODToSSA:units = "None" ;
		NUV_UncertaintyCODToSSA:scale_factor = 0.1 ;
		NUV_UncertaintyCODToSSA:add_offset = 0. ;
		NUV_UncertaintyCODToSSA:Parameter_Type = "Output" ;
		NUV_UncertaintyCODToSSA:Geolocation_Pointer = "Internal geolocation arrays" ;
		NUV_UncertaintyCODToSSA:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		NUV_UncertaintyCODToSSA:_ChunkSizes = 32, 32, 2 ;
		NUV_UncertaintyCODToSSA:_DeflateLevel = 4 ;

    short Quality_flag_Aerosol_Optical_Depth(number_of_lines_7x7, number_of_pixels_7x7) ;
		Quality_flag_Aerosol_Optical_Depth:valid_range = 0s, 3000s ;
		Quality_flag_Aerosol_Optical_Depth:_FillValue = -9999s ;
		Quality_flag_Aerosol_Optical_Depth:long_name = "Land=0 Ocean,0,1,2,3" ;
		Quality_flag_Aerosol_Optical_Depth:units = "None" ;
		Quality_flag_Aerosol_Optical_Depth:scale_factor = 0.001 ;
		Quality_flag_Aerosol_Optical_Depth:add_offset = 0. ;
		Quality_flag_Aerosol_Optical_Depth:Parameter_Type = "Output" ;
		Quality_flag_Aerosol_Optical_Depth:Geolocation_Pointer = "Internal geolocation arrays" ;
		Quality_flag_Aerosol_Optical_Depth:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		Quality_flag_Aerosol_Optical_Depth:_ChunkSizes = 32, 32 ;
		Quality_flag_Aerosol_Optical_Depth:_DeflateLevel = 4 ;
                
    short Quality_flag_SingleScattAlbedo(number_of_lines_7x7, number_of_pixels_7x7) ;
		Quality_flag_SingleScattAlbedo:valid_range = 0s, 3000s ;
		Quality_flag_SingleScattAlbedo:_FillValue = -9999s ;
		Quality_flag_SingleScattAlbedo:long_name = "Quality_flag_SingleScattAlbedo 0,1,2,3" ;
		Quality_flag_SingleScattAlbedo:units = "None" ;
		Quality_flag_SingleScattAlbedo:scale_factor = 0.001 ;
		Quality_flag_SingleScattAlbedo:add_offset = 0. ;
		Quality_flag_SingleScattAlbedo:Parameter_Type = "Output" ;
		Quality_flag_SingleScattAlbedo:Geolocation_Pointer = "Internal geolocation arrays" ;
		Quality_flag_SingleScattAlbedo:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
		Quality_flag_SingleScattAlbedo:_ChunkSizes = 32, 32 ;
		Quality_flag_SingleScattAlbedo:_DeflateLevel = 4 ;

    data:
    } // group geophysical_data
}
