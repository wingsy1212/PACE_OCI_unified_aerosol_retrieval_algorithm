netcdf VNPAERDT {
dimensions:
	number_of_lines_10x10 = UNLIMITED ; //   but varies
	number_of_pixels_10x10 = 135 ;
	number_of_lines_1x1 = UNLIMITED ; //  
	number_of_pixels_1x1 = 2700 ;
	Wavelength_Used_Land_1 = 3 ;
	Wavelength_Used_Land_2 = 4 ;	
	Wavelength_Used_Ocean = 7 ;
	Solution_Index = 9 ;
	Quality_Flag_Num = 2 ;

// global attributes:
        :Conventions = "CF-1.6";
        :format_version = 1; 
        :instrument = "MODIS";
        :platform = "Terra OR AQUA";
        :title = "MODIS"; // look this up
        :processing_level = "L2";
        :processing_version = "v1.0.4";
        :cdm_data_type = "swath";
        :creator_name = "NASA ABI Atmosphere SIPS, Space Science and Engineering Center, University of Wisconsin-Madison";
        :creator_email = "sips.support@ssec.wisc.edu";
        :creator_url = "http://sips.ssec.wisc.edu/";
        :institution = "NASA ABI Atmosphere SIPS";
        :project = "NASA ABI Atmosphere Discipline";
        :publisher_name = "NASA ABI Atmosphere SIPS, Space Science and Engineering Center, University of Wisconsin-Madison";
        :publisher_email = "sips.support@ssec.wisc.edu";
        :publisher_url = "http://sips.ssec.wisc.edu/";
        :keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords";
        :license = "http://science.nasa.gov/earth-science/earth-science-data/data-information-policy/";
        :stdname_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention";
        :naming_authority = "gov.nasa.gsfc.sci.atmos";
        :history = "";
        :source = "";

group: geolocation_data {
    variables:
	float longitude(number_of_lines_10x10, number_of_pixels_10x10) ;
		longitude:valid_range = -180.f, 180.f ;
		longitude:_FillValue = -999.f ;
		longitude:long_name = "Geodetic Longitude" ;
		longitude:units = "degree_east" ;
		longitude:scale_factor = 1. ;
		longitude:add_offset = 0. ;
		longitude:Parameter_Type = "Terra or Aqua Input" ;
		longitude:Geolocation_Pointer = "Geolocation data not applicable" ;
		longitude:_CoordinateAxisType = "Lon" ;
	float latitude(number_of_lines_10x10, number_of_pixels_10x10) ;
		latitude:valid_range = -90.f, 90.f ;
		latitude:_FillValue = -999.f ;
		latitude:long_name = "Geodetic Latitude" ;
		latitude:units = "degree_north" ;
		latitude:scale_factor = 1. ;
		latitude:add_offset = 0. ;
		latitude:Parameter_Type = "Terra or Aqua Input" ;
		latitude:Geolocation_Pointer = "Geolocation data not applicable" ;
		latitude:_CoordinateAxisType = "Lat" ;
	short solar_zenith_angle(number_of_lines_10x10, number_of_pixels_10x10) ;
		solar_zenith_angle:valid_range = 0s, 18000s ;
		solar_zenith_angle:_FillValue = -9999s ;
		solar_zenith_angle:long_name = "Solar Zenith Angle, Cell to Sun" ;
		solar_zenith_angle:units = "degree" ;
		solar_zenith_angle:scale_factor = 0.01 ;
		solar_zenith_angle:add_offset = 0. ;
		solar_zenith_angle:Parameter_Type = "Terra or Aqua Input" ;
		solar_zenith_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		solar_zenith_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short solar_azimuth_angle(number_of_lines_10x10, number_of_pixels_10x10) ;
		solar_azimuth_angle:valid_range = -18000s, 18000s ;
		solar_azimuth_angle:_FillValue = -9999s ;
		solar_azimuth_angle:long_name = "Solar Azimuth Angle, Cell to Sun" ;
		solar_azimuth_angle:units = "degree" ;
		solar_azimuth_angle:scale_factor = 0.01 ;
		solar_azimuth_angle:add_offset = 0. ;
		solar_azimuth_angle:Parameter_Type = "Terra or Aqua Input" ;
		solar_azimuth_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		solar_azimuth_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short sensor_zenith_angle(number_of_lines_10x10, number_of_pixels_10x10) ;
		sensor_zenith_angle:valid_range = 0s, 18000s ;
		sensor_zenith_angle:_FillValue = -9999s ;
		sensor_zenith_angle:long_name = "Sensor Zenith Angle, Cell to Sensor" ;
		sensor_zenith_angle:units = "degree" ;
		sensor_zenith_angle:scale_factor = 0.01 ;
		sensor_zenith_angle:add_offset = 0. ;
		sensor_zenith_angle:Parameter_Type = "Terra or Aqua Input" ;
		sensor_zenith_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		sensor_zenith_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short sensor_azimuth_angle(number_of_lines_10x10, number_of_pixels_10x10) ;
		sensor_azimuth_angle:valid_range = -18000s, 18000s ;
		sensor_azimuth_angle:_FillValue = -9999s ;
		sensor_azimuth_angle:long_name = "Sensor Azimuth Angle, Cell to Sensor" ;
		sensor_azimuth_angle:units = "degree" ;
		sensor_azimuth_angle:scale_factor = 0.01 ;
		sensor_azimuth_angle:add_offset = 0. ;
		sensor_azimuth_angle:Parameter_Type = "Terra or Aqua Input" ;
		sensor_azimuth_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		sensor_azimuth_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Scattering_Angle(number_of_lines_10x10, number_of_pixels_10x10) ;
		Scattering_Angle:valid_range = 0s, 18000s ;
		Scattering_Angle:_FillValue = -9999s ;
		Scattering_Angle:long_name = "Scattering Angle" ;
		Scattering_Angle:units = "Degrees" ;
		Scattering_Angle:scale_factor = 0.01 ;
		Scattering_Angle:add_offset = 0. ;
		Scattering_Angle:Parameter_Type = "Output" ;
		Scattering_Angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		Scattering_Angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Glint_Angle(number_of_lines_10x10, number_of_pixels_10x10) ;
                Glint_Angle:valid_range = 0s, 18000s ;
                Glint_Angle:_FillValue = -9999s ;
                Glint_Angle:long_name = "Glint Angle" ;
                Glint_Angle:units = "Degrees" ;
                Glint_Angle:scale_factor = 0.01 ;
                Glint_Angle:add_offset = 0. ;
                Glint_Angle:Parameter_Type = "Output" ;
                Glint_Angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		Glint_Angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
    data:
    } // group geolocation_data

group: geophysical_data {
    variables:
	short Land_Sea_Flag(number_of_lines_10x10, number_of_pixels_10x10) ;
		Land_Sea_Flag:valid_range = 0s, 1s ;
		Land_Sea_Flag:_FillValue = -9999s ;
		Land_Sea_Flag:long_name = "Land_Sea_Flag(based on MOD03 Landsea mask 0 = Ocean, 1 = Land and ephemeral water 2 = Coastal)" ;
		Land_Sea_Flag:units = "None" ;
		Land_Sea_Flag:scale_factor = 1. ;
		Land_Sea_Flag:add_offset = 0. ;
		Land_Sea_Flag:Parameter_Type = "Output" ;
		Land_Sea_Flag:Geolocation_Pointer = "Internal geolocation arrays" ;
		Land_Sea_Flag:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Aerosol_Cldmask_Land_Ocean(number_of_lines_1x1, number_of_pixels_1x1) ;
		Aerosol_Cldmask_Land_Ocean:valid_range = 0s, 1s ;
		Aerosol_Cldmask_Land_Ocean:_FillValue = -9999s ;
		Aerosol_Cldmask_Land_Ocean:long_name = "Aerosol Cloud Mask at Native resolution  0 = Cloud 1 = Clear" ;
		Aerosol_Cldmask_Land_Ocean:units = "None" ;
		Aerosol_Cldmask_Land_Ocean:scale_factor = 1. ;
		Aerosol_Cldmask_Land_Ocean:add_offset = 0. ;
		Aerosol_Cldmask_Land_Ocean:Parameter_Type = "Output" ;
		Aerosol_Cldmask_Land_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
	short Cloud_Pixel_Distance_Land_Ocean(number_of_lines_1x1, number_of_pixels_1x1) ;
		Cloud_Pixel_Distance_Land_Ocean:valid_range = 0s, 60s ;
		Cloud_Pixel_Distance_Land_Ocean:_FillValue = -9999s ;
		Cloud_Pixel_Distance_Land_Ocean:long_name = "Distance (number of pixels) to nearest pixel identified as cloudy (Native resolution)" ;
		Cloud_Pixel_Distance_Land_Ocean:units = "Number of Pixels" ;
		Cloud_Pixel_Distance_Land_Ocean:scale_factor = 1. ;
		Cloud_Pixel_Distance_Land_Ocean:add_offset = 0. ;
		Cloud_Pixel_Distance_Land_Ocean:Parameter_Type = "Output" ;
		Cloud_Pixel_Distance_Land_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Cloud_Pixel_Distance_Land_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Average_Cloud_Pixel_Distance_Land_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Average_Cloud_Pixel_Distance_Land_Ocean:valid_range = 0s, 60s ;
		Average_Cloud_Pixel_Distance_Land_Ocean:_FillValue = -9999s ;
		Average_Cloud_Pixel_Distance_Land_Ocean:long_name = "Average Distance (number of pixels) to nearest pixel identified as cloudy from each clear pixel used for Aerosol Retrieval in 10 km retrieval box" ; 
		Average_Cloud_Pixel_Distance_Land_Ocean:units = "Number of Pixels" ;
		Average_Cloud_Pixel_Distance_Land_Ocean:scale_factor = 1. ;
		Average_Cloud_Pixel_Distance_Land_Ocean:add_offset = 0. ;
		Average_Cloud_Pixel_Distance_Land_Ocean:Parameter_Type = "Output" ;
		Average_Cloud_Pixel_Distance_Land_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Average_Cloud_Pixel_Distance_Land_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Land_Ocean_Quality_Flag(number_of_lines_10x10, number_of_pixels_10x10) ;
		Land_Ocean_Quality_Flag:valid_range = 0s, 3s ;
		Land_Ocean_Quality_Flag:_FillValue = -9999s ;
		Land_Ocean_Quality_Flag:long_name = "Quality flag for land and ocean aerosol retrievals 0 = Bad  1 = Marginal 2 = Good 3 = Very Good)" ;
		Land_Ocean_Quality_Flag:units = "None" ;
		Land_Ocean_Quality_Flag:scale_factor = 1. ;
		Land_Ocean_Quality_Flag:add_offset = 0. ;
		Land_Ocean_Quality_Flag:Parameter_Type = "Output" ;
		Land_Ocean_Quality_Flag:Geolocation_Pointer = "Internal geolocation arrays" ;
		Land_Ocean_Quality_Flag:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Optical_Depth_Land_And_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Optical_Depth_Land_And_Ocean:valid_range = -100s, 5000s ;
		Optical_Depth_Land_And_Ocean:_FillValue = -9999s ;
		Optical_Depth_Land_And_Ocean:long_name = "AOT at 0.55 micron for both ocean (Average) (Quality flag = 1, 2, 3) and land (corrected) (Quality flag = 3)" ;
		Optical_Depth_Land_And_Ocean:units = "None" ;
		Optical_Depth_Land_And_Ocean:scale_factor = 0.001 ;
		Optical_Depth_Land_And_Ocean:add_offset = 0. ;
		Optical_Depth_Land_And_Ocean:Parameter_Type = "Output" ;
		Optical_Depth_Land_And_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Land_And_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Image_Optical_Depth_Land_And_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Image_Optical_Depth_Land_And_Ocean:valid_range = -100s, 5000s ;
		Image_Optical_Depth_Land_And_Ocean:_FillValue = -9999s ;
		Image_Optical_Depth_Land_And_Ocean:long_name = "AOT at 0.55 micron for both ocean (Average) and land (corrected) with all quality data (Quality flag = 0, 1, 2, 3)" ;
		Image_Optical_Depth_Land_And_Ocean:units = "None" ;
		Image_Optical_Depth_Land_And_Ocean:scale_factor = 0.001 ;
		Image_Optical_Depth_Land_And_Ocean:add_offset = 0. ;
		Image_Optical_Depth_Land_And_Ocean:Parameter_Type = "Output" ;
		Image_Optical_Depth_Land_And_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Image_Optical_Depth_Land_And_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Aerosol_Type_Land(number_of_lines_10x10, number_of_pixels_10x10) ;
		Aerosol_Type_Land:valid_range = 0s, 4s ;
		Aerosol_Type_Land:_FillValue = -9999s ;
		Aerosol_Type_Land:long_name = "Aerosol Type: 1 = Continental, 2 = Moderate Absorption Fine, 3 = Strong Absorption Fine, 4 = Weak Absorption Fine, 5 = Dust Coarse" ;
		Aerosol_Type_Land:units = "None" ;
		Aerosol_Type_Land:scale_factor = 1. ;
		Aerosol_Type_Land:add_offset = 0. ;
		Aerosol_Type_Land:Parameter_Type = "Output" ;
		Aerosol_Type_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Aerosol_Type_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Fitting_Error_Land(number_of_lines_10x10, number_of_pixels_10x10) ;
		Fitting_Error_Land:valid_range = 0s, 1000s ;
		Fitting_Error_Land:_FillValue = -9999s ;
		Fitting_Error_Land:long_name = "Spectral Fitting error for inversion over land" ;
		Fitting_Error_Land:units = "None" ;
		Fitting_Error_Land:scale_factor = 0.001 ;
		Fitting_Error_Land:add_offset = 0. ;
		Fitting_Error_Land:Parameter_Type = "Output" ;
		Fitting_Error_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Fitting_Error_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Surface_Reflectance_Land(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Land_1) ;
		Surface_Reflectance_Land:valid_range = 0s, 1000s ;
		Surface_Reflectance_Land:_FillValue = -9999s ;
		Surface_Reflectance_Land:long_name = "Estimated Surface Reflectance at 0.48, 0.67, 2.25 microns" ;
		Surface_Reflectance_Land:units = "None" ;
		Surface_Reflectance_Land:scale_factor = 0.001 ;
		Surface_Reflectance_Land:add_offset = 0. ;
		Surface_Reflectance_Land:Parameter_Type = "Output" ;
		Surface_Reflectance_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Surface_Reflectance_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude " ;
	short Corrected_Optical_Depth_Land(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Land_2) ;
		Corrected_Optical_Depth_Land:valid_range = -100s, 5000s ;
		Corrected_Optical_Depth_Land:_FillValue = -9999s ;
		Corrected_Optical_Depth_Land:long_name = "Retrieved AOT at 0.48, 0.55, 0.67, 2.25 microns" ;
		Corrected_Optical_Depth_Land:units = "None" ;
		Corrected_Optical_Depth_Land:scale_factor = 0.001 ;
		Corrected_Optical_Depth_Land:add_offset = 0. ;
		Corrected_Optical_Depth_Land:Parameter_Type = "Output" ;
		Corrected_Optical_Depth_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Corrected_Optical_Depth_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude " ;
	short Optical_Depth_Ratio_Small_Land(number_of_lines_10x10, number_of_pixels_10x10) ;
		Optical_Depth_Ratio_Small_Land:valid_range = 0s, 1000s ;
		Optical_Depth_Ratio_Small_Land:_FillValue = -9999s ;
		Optical_Depth_Ratio_Small_Land:long_name = "Fraction of AOT contributed by fine dominated model" ;
		Optical_Depth_Ratio_Small_Land:units = "None" ;
		Optical_Depth_Ratio_Small_Land:scale_factor = 0.001 ;
		Optical_Depth_Ratio_Small_Land:add_offset = 0. ;
		Optical_Depth_Ratio_Small_Land:Parameter_Type = "Output" ;
		Optical_Depth_Ratio_Small_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Ratio_Small_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Number_Pixels_Used_Land(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Land_1) ;
		Number_Pixels_Used_Land:valid_range = 1s, 400s ;
		Number_Pixels_Used_Land:_FillValue = -9999s ;
		Number_Pixels_Used_Land:long_name = "Number of pixels used for land retrieval at 0.48,0.67and 2.25 micron " ;
		Number_Pixels_Used_Land:units = "None" ;
		Number_Pixels_Used_Land:scale_factor = 1. ;
		Number_Pixels_Used_Land:add_offset = 0. ;
		Number_Pixels_Used_Land:Parameter_Type = "Output" ;
		Number_Pixels_Used_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Number_Pixels_Used_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Mean_Reflectance_Land(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Land_1) ;
		Mean_Reflectance_Land:valid_range = 0s, 10000s ;
		Mean_Reflectance_Land:_FillValue = -9999s ;
		Mean_Reflectance_Land:long_name = "Mean reflectance of pixels used for land retrieval at 0.48,0.67,2.25  microns " ;
		Mean_Reflectance_Land:units = "None" ;
		Mean_Reflectance_Land:scale_factor = 0.0001 ;
		Mean_Reflectance_Land:add_offset = 0. ;
		Mean_Reflectance_Land:Parameter_Type = "Output" ;
		Mean_Reflectance_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mean_Reflectance_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short STD_Reflectance_Land(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Land_1) ;
		STD_Reflectance_Land:valid_range = 0s, 20000s ;
		STD_Reflectance_Land:_FillValue = -9999s ;
		STD_Reflectance_Land:long_name = "Standard deviation of reflectance of pixels used for land retrieval used for land retrieval at 0.48,0.67,2.25  microns " ;
		STD_Reflectance_Land:units = "None" ;
		STD_Reflectance_Land:scale_factor = 0.0001 ;
		STD_Reflectance_Land:add_offset = 0. ;
		STD_Reflectance_Land:Parameter_Type = "Output" ;
		STD_Reflectance_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		STD_Reflectance_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	float Mass_Concentration_Land(number_of_lines_10x10, number_of_pixels_10x10) ;
		Mass_Concentration_Land:valid_range = 0.f, 1000.f ;
		Mass_Concentration_Land:_FillValue = -999.f ;
		Mass_Concentration_Land:long_name = "Estimated Column Mass(per area) using assumed mass extinction efficiency" ;
		Mass_Concentration_Land:units = "1.0e-6g/cm^2" ;
		Mass_Concentration_Land:scale_factor = 1. ;
		Mass_Concentration_Land:add_offset = 0. ;
		Mass_Concentration_Land:Parameter_Type = "Output" ;
		Mass_Concentration_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mass_Concentration_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Aerosol_Cloud_Fraction_Land(number_of_lines_10x10, number_of_pixels_10x10) ;
		Aerosol_Cloud_Fraction_Land:valid_range = 0s, 1000s ;
		Aerosol_Cloud_Fraction_Land:_FillValue = -9999s ;
		Aerosol_Cloud_Fraction_Land:long_name = "Cloud fraction from Land aerosol cloud mask from retrieved and overcast pixels not including cirrus mask" ;
		Aerosol_Cloud_Fraction_Land:units = "None" ;
		Aerosol_Cloud_Fraction_Land:scale_factor = 0.001 ;
		Aerosol_Cloud_Fraction_Land:add_offset = 0. ;
		Aerosol_Cloud_Fraction_Land:Parameter_Type = "Output" ;
		Aerosol_Cloud_Fraction_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Aerosol_Cloud_Fraction_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Effective_Optical_Depth_Average_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Ocean) ;
		Effective_Optical_Depth_Average_Ocean:valid_range = -100s, 5000s ;
		Effective_Optical_Depth_Average_Ocean:_FillValue = -9999s ;
		Effective_Optical_Depth_Average_Ocean:long_name = "Retrieved AOT for  average  solution at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Effective_Optical_Depth_Average_Ocean:units = "None" ;
		Effective_Optical_Depth_Average_Ocean:scale_factor = 0.001 ;
		Effective_Optical_Depth_Average_Ocean:add_offset = 0. ;
		Effective_Optical_Depth_Average_Ocean:Parameter_Type = "Output" ;
		Effective_Optical_Depth_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Effective_Optical_Depth_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Optical_Depth_Small_Average_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Ocean) ;
		Optical_Depth_Small_Average_Ocean:valid_range = -100s, 5000s ;
		Optical_Depth_Small_Average_Ocean:_FillValue = -9999s ;
		Optical_Depth_Small_Average_Ocean:long_name = "Retrieved optical thickness for fine mode (Average solution) for 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Optical_Depth_Small_Average_Ocean:units = "None" ;
		Optical_Depth_Small_Average_Ocean:scale_factor = 0.001 ;
		Optical_Depth_Small_Average_Ocean:add_offset = 0. ;
		Optical_Depth_Small_Average_Ocean:Parameter_Type = "Output" ;
		Optical_Depth_Small_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Small_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Optical_Depth_Large_Average_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Ocean) ;
		Optical_Depth_Large_Average_Ocean:valid_range = -100s, 5000s ;
		Optical_Depth_Large_Average_Ocean:_FillValue = -9999s ;
		Optical_Depth_Large_Average_Ocean:long_name = "Retrieved AOT of large mode for  average  solution at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Optical_Depth_Large_Average_Ocean:units = "None" ;
		Optical_Depth_Large_Average_Ocean:scale_factor = 0.001 ;
		Optical_Depth_Large_Average_Ocean:add_offset = 0. ;
		Optical_Depth_Large_Average_Ocean:Parameter_Type = "Output" ;
		Optical_Depth_Large_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Large_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	float Mass_Concentration_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Mass_Concentration_Ocean:valid_range = 0.f, 1000.f ;
		Mass_Concentration_Ocean:_FillValue = -999.f ;
		Mass_Concentration_Ocean:long_name = "Estimated Column Mass (per area) using assumed mass extinction coefficients" ;
		Mass_Concentration_Ocean:units = "1.0e-6g/cm^2" ;
		Mass_Concentration_Ocean:scale_factor = 1. ;
		Mass_Concentration_Ocean:add_offset = 0. ;
		Mass_Concentration_Ocean:Parameter_Type = "Output" ;
		Mass_Concentration_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mass_Concentration_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Aerosol_Cloud_Fraction_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Aerosol_Cloud_Fraction_Ocean:valid_range = 0s, 1000s ;
		Aerosol_Cloud_Fraction_Ocean:_FillValue = -9999s ;
		Aerosol_Cloud_Fraction_Ocean:long_name = "Cloud fraction from Ocean aerosol cloud mask from retrieved and overcast pixels not including cirrus mask" ;
		Aerosol_Cloud_Fraction_Ocean:units = "None" ;
		Aerosol_Cloud_Fraction_Ocean:scale_factor = 0.001 ;
		Aerosol_Cloud_Fraction_Ocean:add_offset = 0. ;
		Aerosol_Cloud_Fraction_Ocean:Parameter_Type = "Output" ;
		Aerosol_Cloud_Fraction_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Aerosol_Cloud_Fraction_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Effective_Radius_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Effective_Radius_Ocean:valid_range = 0s, 5000s ;
		Effective_Radius_Ocean:_FillValue = -9999s ;
		Effective_Radius_Ocean:long_name = "Effective_Radius at 0.55 microns" ;
		Effective_Radius_Ocean:units = "micron" ;
		Effective_Radius_Ocean:scale_factor = 0.001 ;
		Effective_Radius_Ocean:add_offset = 0. ;
		Effective_Radius_Ocean:Parameter_Type = "Output" ;
		Effective_Radius_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Effective_Radius_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	float PSML003_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		PSML003_Ocean:valid_range = 0.f, 9.9999998e+10f ;
		PSML003_Ocean:_FillValue = -999.f ;
		PSML003_Ocean:long_name = "Inferred column number concentration (number per area) of particles larger than 0.03 micron " ;
		PSML003_Ocean:units = "Particles/cm^2" ;
		PSML003_Ocean:scale_factor = 1. ;
		PSML003_Ocean:add_offset = 0. ;
		PSML003_Ocean:Parameter_Type = "Output" ;
		PSML003_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		PSML003_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Asymmetry_Factor_Average_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Ocean) ;
		Asymmetry_Factor_Average_Ocean:valid_range = 0s, 3000s ;
		Asymmetry_Factor_Average_Ocean:_FillValue = -9999s ;
		Asymmetry_Factor_Average_Ocean:long_name = "Inferred Asymmetry_Factor for  average  solution at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Asymmetry_Factor_Average_Ocean:units = "None" ;
		Asymmetry_Factor_Average_Ocean:scale_factor = 0.001 ;
		Asymmetry_Factor_Average_Ocean:add_offset = 0. ;
		Asymmetry_Factor_Average_Ocean:Parameter_Type = "Output" ;
		Asymmetry_Factor_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Asymmetry_Factor_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Backscattering_Ratio_Average_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Ocean) ;
		Backscattering_Ratio_Average_Ocean:valid_range = 0s, 3000s ;
		Backscattering_Ratio_Average_Ocean:_FillValue = -9999s ;
		Backscattering_Ratio_Average_Ocean:long_name = "Inferred Backscattering_Ratio for  average  solution at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Backscattering_Ratio_Average_Ocean:units = "None" ;
		Backscattering_Ratio_Average_Ocean:scale_factor = 0.001 ;
		Backscattering_Ratio_Average_Ocean:add_offset = 0. ;
		Backscattering_Ratio_Average_Ocean:Parameter_Type = "Output" ;
		Backscattering_Ratio_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Backscattering_Ratio_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Angstrom_Exponent_1_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Angstrom_Exponent_1_Ocean:valid_range = -1000s, 5000s ;
		Angstrom_Exponent_1_Ocean:_FillValue = -9999s ;
		Angstrom_Exponent_1_Ocean:long_name = "Calculated Angstrom Exponent for 0.55 vs 0.86 micron  for Average Solution" ;
		Angstrom_Exponent_1_Ocean:units = "None" ;
		Angstrom_Exponent_1_Ocean:scale_factor = 0.001 ;
		Angstrom_Exponent_1_Ocean:add_offset = 0. ;
		Angstrom_Exponent_1_Ocean:Parameter_Type = "Output" ;
		Angstrom_Exponent_1_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Angstrom_Exponent_1_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Angstrom_Exponent_2_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Angstrom_Exponent_2_Ocean:valid_range = -1000s, 5000s ;
		Angstrom_Exponent_2_Ocean:_FillValue = -9999s ;
		Angstrom_Exponent_2_Ocean:long_name = "Calculated Angstrom Exponent for 0.86 vs 2.13 micron for Average Solution" ;
		Angstrom_Exponent_2_Ocean:units = "None" ;
		Angstrom_Exponent_2_Ocean:scale_factor = 0.001 ;
		Angstrom_Exponent_2_Ocean:add_offset = 0. ;
		Angstrom_Exponent_2_Ocean:Parameter_Type = "Output" ;
		Angstrom_Exponent_2_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Angstrom_Exponent_2_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Least_Squares_Error_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Least_Squares_Error_Ocean:valid_range = 0s, 1000s ;
		Least_Squares_Error_Ocean:_FillValue = -9999s ;
		Least_Squares_Error_Ocean:long_name = "Residual of least squares fitting for inversion over ocean" ;
		Least_Squares_Error_Ocean:units = "None" ;
		Least_Squares_Error_Ocean:scale_factor = 0.001 ;
		Least_Squares_Error_Ocean:add_offset = 0. ;
		Least_Squares_Error_Ocean:Parameter_Type = "Output" ;
		Least_Squares_Error_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Least_Squares_Error_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Optical_Depth_Ratio_Small_Ocean_0p55micron(number_of_lines_10x10, number_of_pixels_10x10) ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:valid_range = 0s, 1000s ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:_FillValue = -9999s ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:long_name = "Fraction of AOT (at 0.55 micron) contributed by fine mode for average solution" ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:units = "None" ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:scale_factor = 0.001 ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:add_offset = 0. ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:Parameter_Type = "Output" ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Optical_Depth_By_Models_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Solution_Index) ;
		Optical_Depth_By_Models_Ocean:valid_range = -100s, 5000s ;
		Optical_Depth_By_Models_Ocean:_FillValue = -9999s ;
		Optical_Depth_By_Models_Ocean:long_name = "Retrieved AOT (at 0.55 micron) partioned by mode index (for Best solution)" ;
		Optical_Depth_By_Models_Ocean:units = "None" ;
		Optical_Depth_By_Models_Ocean:scale_factor = 0.001 ;
		Optical_Depth_By_Models_Ocean:add_offset = 0. ;
		Optical_Depth_By_Models_Ocean:Parameter_Type = "Output" ;
		Optical_Depth_By_Models_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_By_Models_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Number_Pixels_Used_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Ocean) ;
		Number_Pixels_Used_Ocean:valid_range = 1s, 400s ;
		Number_Pixels_Used_Ocean:_FillValue = -9999s ;
		Number_Pixels_Used_Ocean:long_name = "Number of pixels used for ocean retrieval at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 micron)" ;
		Number_Pixels_Used_Ocean:units = "None" ;
		Number_Pixels_Used_Ocean:scale_factor = 1. ;
		Number_Pixels_Used_Ocean:add_offset = 0. ;
		Number_Pixels_Used_Ocean:Parameter_Type = "Output" ;
		Number_Pixels_Used_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Number_Pixels_Used_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Mean_Reflectance_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Ocean) ;
		Mean_Reflectance_Ocean:valid_range = 0s, 10000s ;
		Mean_Reflectance_Ocean:_FillValue = -9999s ;
		Mean_Reflectance_Ocean:long_name = "Mean reflectance of pixels used for ocean retrieval at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 micron " ;
		Mean_Reflectance_Ocean:units = "None" ;
		Mean_Reflectance_Ocean:scale_factor = 0.0001 ;
		Mean_Reflectance_Ocean:add_offset = 0. ;
		Mean_Reflectance_Ocean:Parameter_Type = "Output" ;
		Mean_Reflectance_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mean_Reflectance_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short STD_Reflectance_Ocean(number_of_lines_10x10, number_of_pixels_10x10, Wavelength_Used_Ocean) ;
		STD_Reflectance_Ocean:valid_range = 0s, 20000s ;
		STD_Reflectance_Ocean:_FillValue = -9999s ;
		STD_Reflectance_Ocean:long_name = "Standard deviation of reflectance of pixels used for ocean retrieval at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns )" ;
		STD_Reflectance_Ocean:units = "None" ;
		STD_Reflectance_Ocean:scale_factor = 0.0001 ;
		STD_Reflectance_Ocean:add_offset = 0. ;
		STD_Reflectance_Ocean:Parameter_Type = "Output" ;
		STD_Reflectance_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		STD_Reflectance_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Wind_Speed_Ncep_Ocean(number_of_lines_10x10, number_of_pixels_10x10) ;
		Wind_Speed_Ncep_Ocean:valid_range = 0s, 8000s ;
		Wind_Speed_Ncep_Ocean:_FillValue = -9999s ;
		Wind_Speed_Ncep_Ocean:long_name = "Wind Speed based on NCEP reanalysis for Ocean" ;
		Wind_Speed_Ncep_Ocean:units = "Meters/sec" ;
		Wind_Speed_Ncep_Ocean:scale_factor = 0.01 ;
		Wind_Speed_Ncep_Ocean:add_offset = 0. ;
		Wind_Speed_Ncep_Ocean:Parameter_Type = "Output" ;
		Wind_Speed_Ncep_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Wind_Speed_Ncep_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Topographic_Altitude_Land(number_of_lines_10x10, number_of_pixels_10x10) ;
		Topographic_Altitude_Land:valid_range = 0s, 1000s ;
		Topographic_Altitude_Land:_FillValue = -9999s ;
		Topographic_Altitude_Land:long_name = "Averaged topographic altitude (in km) for Land" ;
		Topographic_Altitude_Land:units = "KM" ;
		Topographic_Altitude_Land:scale_factor = 0.01 ;
		Topographic_Altitude_Land:add_offset = 0. ;
		Topographic_Altitude_Land:Parameter_Type = "Output" ;
		Topographic_Altitude_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Topographic_Altitude_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
	short Error_Flag_Land_And_Ocean(number_of_lines_10x10, number_of_pixels_10x10,Quality_Flag_Num) ;
		Error_Flag_Land_And_Ocean:valid_range = 1s, 26s ;
                Error_Flag_Land_And_Ocean:_FillValue = -9999s ;
                Error_Flag_Land_And_Ocean:long_name = "Error code 1-26. Layer 1 ocean, Layer 2 land. Ask for Documentation" ;
                Error_Flag_Land_And_Ocean:units = "None" ;
                Error_Flag_Land_And_Ocean:scale_factor = 1.0 ;
                Error_Flag_Land_And_Ocean:add_offset = 0. ;
                Error_Flag_Land_And_Ocean:Parameter_Type = "Output" ;
                Error_Flag_Land_And_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Error_Flag_Land_And_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
    data:
    } // group geophysical_data
}
