netcdf AERDT_L2_OCI {
dimensions:
	number_of_lines = UNLIMITED ; // e.g. 3232
	pixels_per_line = 1272 ;
	Wavelength_Used_UV1 = 2 ;
// global attributes:
        :Conventions = "CF-1.8 ACDD-1.3";
        :format_version = 1;
        :instrument = "OCI";
        :platform = "PACE";  // Suomi-NPP or NOAA-20
        :processing_level = "L2";
        :processing_version = "";
        :cdm_data_type = "swath";
        :creator_name = "NASA/GSFC/OBPG";
        :creator_email = "data@oceancolor.gsfc.nasa.gov";
        :creator_url = "https://oceandata.sci.gsfc.nasa.gov";
        :institution = "NASA Goddard Space Flight Center, Ocean Biology Processing Group";
        :project = "Ocean Biology Processing Group (NASA/GSFC/OBPG)";
        :publisher_name = "NASA/GSFC/OBPG";
        :publisher_email = "data@oceancolor.gsfc.nasa.gov";
        :publisher_url = "https://oceandata.sci.gsfc.nasa.gov";
        :keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords";
        :license = "https://science.nasa.gov/earth-science/earth-science-data/data-information-policy/";
        :stdname_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention";
        :naming_authority = "gov.nasa.gsfc.sci.oceandata";
        :title = "PACE OCI Level-2 Data UAA 1x1";

group: processing_control {
        // No dimensions or variables needed
        :software_name = "OCI Unified Aerosol Algorithm (UAA)";
        :software_version = "3.0.0";
        :config_file = "";
    } // group processing_control

group: geolocation_data {
    variables:
	float Longitude_1km(number_of_lines, pixels_per_line) ;
		Longitude_1km:valid_range = -180.f, 180.f ;
		Longitude_1km:_FillValue = -999.f ;
		Longitude_1km:long_name = "Geodetic Longitude_1km" ;
		Longitude_1km:units = "degree_east" ;
		Longitude_1km:_CoordinateAxisType = "Lon" ;
		Longitude_1km:_ChunkSizes = 128, 128 ;
		Longitude_1km:_DeflateLevel = 4 ;

	float Latitude_1km(number_of_lines, pixels_per_line) ;
		Latitude_1km:valid_range = -90.f, 90.f ;
		Latitude_1km:_FillValue = -999.f ;
		Latitude_1km:long_name = "Geodetic Latitude_1km" ;
		Latitude_1km:units = "degree_north" ;
		Latitude_1km:_CoordinateAxisType = "Lat" ;
		Latitude_1km:_ChunkSizes = 128, 128 ;
		Latitude_1km:_DeflateLevel = 4 ;


    data:
    } // group geolocation_data
group: geophysical_data {
    variables:


	short NUV_AerosolIndex_1km(number_of_lines, pixels_per_line) ;
		NUV_AerosolIndex_1km:valid_range =  -5000s, 10000s ;
		NUV_AerosolIndex_1km:_FillValue = -9999s ;
		NUV_AerosolIndex_1km:long_name = "NUV Retrieved Aerosol Index (0.354,0.388) Pair at native 1km resolution"  ;
		NUV_AerosolIndex_1km:scale_factor = 0.001 ;
		NUV_AerosolIndex_1km:add_offset = 0. ;
		NUV_AerosolIndex_1km:coordinates = "/geolocation_data/Longitude_1km /geolocation_data/Latitude_1km" ;
		NUV_AerosolIndex_1km:_ChunkSizes = 128, 128 ;
		NUV_AerosolIndex_1km:_DeflateLevel = 4 ;

	short NUV_Residue_1km(number_of_lines, pixels_per_line) ;
		NUV_Residue_1km:valid_range =  -5000s, 10000s ;
		NUV_Residue_1km:_FillValue = -9999s ;
		NUV_Residue_1km:long_name = "NUV Retrieved LER based AI (0.354,0.388) Pair at native 1km resolution"  ;
		NUV_Residue_1km:scale_factor = 0.001 ;
		NUV_Residue_1km:add_offset = 0. ;
		NUV_Residue_1km:coordinates = "/geolocation_data/Longitude_1km /geolocation_data/Latitude_1km" ;
		NUV_Residue_1km:_ChunkSizes = 128, 128 ;
		NUV_Residue_1km:_DeflateLevel = 4 ;

	short NUV_Reflectivity_1km(number_of_lines, pixels_per_line, Wavelength_Used_UV1) ;
		NUV_Reflectivity_1km:valid_range =  0s, 1000s ;
		NUV_Reflectivity_1km:_FillValue = -9999s ;
		NUV_Reflectivity_1km:long_name = "NUV Retrieved LERs for 0.354 and 0.388 micron at native 1km resolution"  ;
		NUV_Reflectivity_1km:scale_factor = 0.001 ;
		NUV_Reflectivity_1km:add_offset = 0. ;
		NUV_Reflectivity_1km:coordinates = "/geolocation_data/Longitude_1km /geolocation_data/Latitude_1km" ;
		NUV_Reflectivity_1km:_ChunkSizes = 128, 128, 2 ;
		NUV_Reflectivity_1km:_DeflateLevel = 4 ;

    data:
    } // group geophysical_data
}
