netcdf AERDT_L2_VIIRS {
dimensions:
	number_of_lines_8x8 = UNLIMITED ; // e.g. 404 but varies
	number_of_pixels_8x8 = 400 ;
	number_of_lines_1x1 = UNLIMITED ; // e.g. 3232
	number_of_pixels_1x1 = 2000;
	Wavelength_Used_Land_1 = 3 ;
	Wavelength_Used_Land_2 = 4 ;
	Wavelength_Used_Land_3 = 7 ;
	Wavelength_Used_Ocean = 7 ;
	Solution_Index = 10 ;
	Quality_Flag_Num = 2 ;

// global attributes:
        :Conventions = "CF-1.6";
        :format_version = 1; 
        :instrument = "VIIRS";
        :platform = "";  // Suomi-NPP or NOAA-20
        :processing_level = "L2";
        :cdm_data_type = "swath";
        :creator_name = "NASA Atmosphere SIPS";
        :creator_email = "sips.support@ssec.wisc.edu";
        :creator_url = "https://sips.ssec.wisc.edu/";
        :institution = "NASA Atmosphere SIPS";
        :project = "NASA Atmosphere Discipline";
        :publisher_name = "NASA Atmosphere SIPS";
        :publisher_email = "sips.support@ssec.wisc.edu";
        :publisher_url = "https://sips.ssec.wisc.edu/";
        :date_created = "";
        :product_name = "";
        :LocalGranuleID = "";
        :ShortName = "AERDT_L2_VIIRS_SNPP";
        :product_version = ""; // if operational
        :identifier_product_doi = ""; // if operational
	:identifier_product_doi_authority = "http://dx.doi.org";
        :ancillary_files = "";
        :l1_version = "";
        :l1_lut_version = "";
        :l1_lut_created = "";
	:DataCenterId = "UWI-MAD/SSEC/ASIPS";
	:creator_institution = "Space Science & Engineering Center, University of Wisconsin - Madison";
	:publisher_institution = "NASA Level-1 and Atmosphere Archive & Distribution System";
        :keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords";
        :license = "https://science.nasa.gov/earth-science/earth-science-data/data-information-policy/";
        :stdname_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention";
        :naming_authority = "gov.nasa.gsfc.sci.atmos";
        :history = "";
        :source = "";
        :title = "SNPP Dark Target Aerosol (AERDT_L2_VIIRS_SNPP)";
        :long_name = "SNPP VIIRS Dark Target Aerosol 6-Min L2 Swath 6 km";
        :processing_version = "";
        :l2_lut_files = "big_v1c1.dat.npp4,big_v2c1.dat.npp4,big_v3c1.dat.npp4,big_v4c1.dat.npp4,small_v1c1.dat.npp4,small_v2c1.dat.npp4,small_v3c1.dat.npp4,small_v4c1.dat.npp4,Ocean_Ext_554_modislike,lookup_land_w0488.npp3,lookup_land_w0551.npp3,lookup_land_w0670.npp3,lookup_land_w2257.npp3,Urban_Table_10km,aerosol_land_map.v3";

group: geolocation_data {
    variables:
	float longitude(number_of_lines_8x8, number_of_pixels_8x8) ;
		longitude:valid_range = -180.f, 180.f ;
		longitude:_FillValue = -999.f ;
		longitude:long_name = "Geodetic Longitude" ;
		longitude:units = "degree_east" ;
		longitude:scale_factor = 1. ;
		longitude:add_offset = 0. ;
		longitude:Parameter_Type = "VIIRS Input" ;
		longitude:Geolocation_Pointer = "Geolocation data not applicable" ;
		longitude:_CoordinateAxisType = "Lon" ;
        longitude:_Storage = "chunked" ;
        longitude:_ChunkSizes = 1, 400 ;
        longitude:_DeflateLevel = 5 ;
        longitude:_Shuffle = "true" ;
	float latitude(number_of_lines_8x8, number_of_pixels_8x8) ;
		latitude:valid_range = -90.f, 90.f ;
		latitude:_FillValue = -999.f ;
		latitude:long_name = "Geodetic Latitude" ;
		latitude:units = "degree_north" ;
		latitude:scale_factor = 1. ;
		latitude:add_offset = 0. ;
		latitude:Parameter_Type = "VIIRS Input" ;
		latitude:Geolocation_Pointer = "Geolocation data not applicable" ;
		latitude:_CoordinateAxisType = "Lat" ;
        latitude:_Storage = "chunked" ;
        latitude:_ChunkSizes = 1, 400 ;
        latitude:_DeflateLevel = 5 ;
        latitude:_Shuffle = "true" ;
	short solar_zenith_angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		solar_zenith_angle:valid_range = 0s, 18000s ;
		solar_zenith_angle:_FillValue = -9999s ;
		solar_zenith_angle:long_name = "Solar Zenith Angle, Cell to Sun" ;
		solar_zenith_angle:units = "degree" ;
		solar_zenith_angle:scale_factor = 0.01 ;
		solar_zenith_angle:add_offset = 0. ;
		solar_zenith_angle:Parameter_Type = "VIIRS Input" ;
		solar_zenith_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		solar_zenith_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        solar_zenith_angle:_Storage = "chunked" ;
        solar_zenith_angle:_ChunkSizes = 1, 400 ;
        solar_zenith_angle:_DeflateLevel = 5 ;
        solar_zenith_angle:_Shuffle = "true" ;
	short solar_azimuth_angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		solar_azimuth_angle:valid_range = -18000s, 18000s ;
		solar_azimuth_angle:_FillValue = -9999s ;
		solar_azimuth_angle:long_name = "Solar Azimuth Angle, Cell to Sun" ;
		solar_azimuth_angle:units = "degree" ;
		solar_azimuth_angle:scale_factor = 0.01 ;
		solar_azimuth_angle:add_offset = 0. ;
		solar_azimuth_angle:Parameter_Type = "VIIRS Input" ;
		solar_azimuth_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		solar_azimuth_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        solar_azimuth_angle:_Storage = "chunked" ;
        solar_azimuth_angle:_ChunkSizes = 1, 400 ;
        solar_azimuth_angle:_DeflateLevel = 5 ;
        solar_azimuth_angle:_Shuffle = "true" ;
	short sensor_zenith_angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		sensor_zenith_angle:valid_range = 0s, 18000s ;
		sensor_zenith_angle:_FillValue = -9999s ;
		sensor_zenith_angle:long_name = "Sensor Zenith Angle, Cell to Sensor" ;
		sensor_zenith_angle:units = "degree" ;
		sensor_zenith_angle:scale_factor = 0.01 ;
		sensor_zenith_angle:add_offset = 0. ;
		sensor_zenith_angle:Parameter_Type = "VIIRS Input" ;
		sensor_zenith_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		sensor_zenith_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        sensor_zenith_angle:_Storage = "chunked" ;
        sensor_zenith_angle:_ChunkSizes = 1, 400 ;
        sensor_zenith_angle:_DeflateLevel = 5 ;
        sensor_zenith_angle:_Shuffle = "true" ;
	short sensor_azimuth_angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		sensor_azimuth_angle:valid_range = -18000s, 18000s ;
		sensor_azimuth_angle:_FillValue = -9999s ;
		sensor_azimuth_angle:long_name = "Sensor Azimuth Angle, Cell to Sensor" ;
		sensor_azimuth_angle:units = "degree" ;
		sensor_azimuth_angle:scale_factor = 0.01 ;
		sensor_azimuth_angle:add_offset = 0. ;
		sensor_azimuth_angle:Parameter_Type = "VIIRS Input" ;
		sensor_azimuth_angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		sensor_azimuth_angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        sensor_azimuth_angle:_Storage = "chunked" ;
        sensor_azimuth_angle:_ChunkSizes = 1, 400 ;
        sensor_azimuth_angle:_DeflateLevel = 5 ;
        sensor_azimuth_angle:_Shuffle = "true" ;
	short Scattering_Angle(number_of_lines_8x8, number_of_pixels_8x8) ;
		Scattering_Angle:valid_range = 0s, 18000s ;
		Scattering_Angle:_FillValue = -9999s ;
		Scattering_Angle:long_name = "Scattering Angle" ;
		Scattering_Angle:units = "Degrees" ;
		Scattering_Angle:scale_factor = 0.01 ;
		Scattering_Angle:add_offset = 0. ;
		Scattering_Angle:Parameter_Type = "Output" ;
		Scattering_Angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		Scattering_Angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Scattering_Angle:_Storage = "chunked" ;
        Scattering_Angle:_ChunkSizes = 1, 400 ;
        Scattering_Angle:_DeflateLevel = 5 ;
        Scattering_Angle:_Shuffle = "true" ;
	short Glint_Angle(number_of_lines_8x8, number_of_pixels_8x8) ;
        Glint_Angle:valid_range = 0s, 18000s ;
        Glint_Angle:_FillValue = -9999s ;
        Glint_Angle:long_name = "Glint Angle" ;
        Glint_Angle:units = "Degrees" ;
        Glint_Angle:scale_factor = 0.01 ;
        Glint_Angle:add_offset = 0. ;
        Glint_Angle:Parameter_Type = "Output" ;
        Glint_Angle:Geolocation_Pointer = "Internal geolocation arrays" ;
		Glint_Angle:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Glint_Angle:_Storage = "chunked" ;
        Glint_Angle:_ChunkSizes = 1, 400 ;
        Glint_Angle:_DeflateLevel = 5 ;
        Glint_Angle:_Shuffle = "true" ;
    data:
    } // group geolocation_data

group: geophysical_data {
    variables:
	short Land_Sea_Flag(number_of_lines_8x8, number_of_pixels_8x8) ;
		Land_Sea_Flag:valid_range = 0s, 1s ;
		Land_Sea_Flag:_FillValue = -9999s ;
		Land_Sea_Flag:long_name = "Land_Sea_Flag(based on MOD03 Landsea mask 0 = Ocean, 1 = Land and ephemeral water 2 = Coastal)" ;
		Land_Sea_Flag:units = "None" ;
		Land_Sea_Flag:scale_factor = 1. ;
		Land_Sea_Flag:add_offset = 0. ;
		Land_Sea_Flag:Parameter_Type = "Output" ;
		Land_Sea_Flag:Geolocation_Pointer = "Internal geolocation arrays" ;
		Land_Sea_Flag:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Land_Sea_Flag:_Storage = "chunked" ;
        Land_Sea_Flag:_ChunkSizes = 1, 400 ;
        Land_Sea_Flag:_DeflateLevel = 5 ;
        Land_Sea_Flag:_Shuffle = "true" ;
	short Aerosol_Cldmask_Land_Ocean(number_of_lines_1x1, number_of_pixels_1x1) ;
		Aerosol_Cldmask_Land_Ocean:valid_range = 0s, 1s ;
		Aerosol_Cldmask_Land_Ocean:_FillValue = -9999s ;
		Aerosol_Cldmask_Land_Ocean:long_name = "Aerosol Cloud Mask 750 meter resolution 0 = Cloud 1 = Clear" ;
		Aerosol_Cldmask_Land_Ocean:units = "None" ;
		Aerosol_Cldmask_Land_Ocean:scale_factor = 1. ;
		Aerosol_Cldmask_Land_Ocean:add_offset = 0. ;
		Aerosol_Cldmask_Land_Ocean:Parameter_Type = "Output" ;
		Aerosol_Cldmask_Land_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
        Aerosol_Cldmask_Land_Ocean:_Storage = "chunked" ;
        Aerosol_Cldmask_Land_Ocean:_ChunkSizes = 1, 400 ;
        Aerosol_Cldmask_Land_Ocean:_DeflateLevel = 5 ;
        Aerosol_Cldmask_Land_Ocean:_Shuffle = "true" ;
	short Cloud_Pixel_Distance_Land_Ocean(number_of_lines_1x1, number_of_pixels_1x1) ;
		Cloud_Pixel_Distance_Land_Ocean:valid_range = 0s, 60s ;
		Cloud_Pixel_Distance_Land_Ocean:_FillValue = -9999s ;
		Cloud_Pixel_Distance_Land_Ocean:long_name = "Distance (number of pixels) to nearest pixel identified as cloudy (750 m resolution)" ;
		Cloud_Pixel_Distance_Land_Ocean:units = "Number of Pixels" ;
		Cloud_Pixel_Distance_Land_Ocean:scale_factor = 1. ;
		Cloud_Pixel_Distance_Land_Ocean:add_offset = 0. ;
		Cloud_Pixel_Distance_Land_Ocean:Parameter_Type = "Output" ;
		Cloud_Pixel_Distance_Land_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Cloud_Pixel_Distance_Land_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Cloud_Pixel_Distance_Land_Ocean:_Storage = "chunked" ;
        Cloud_Pixel_Distance_Land_Ocean:_ChunkSizes = 1, 400 ;
        Cloud_Pixel_Distance_Land_Ocean:_DeflateLevel = 5 ;
        Cloud_Pixel_Distance_Land_Ocean:_Shuffle = "true" ;
	short Average_Cloud_Pixel_Distance_Land_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Average_Cloud_Pixel_Distance_Land_Ocean:valid_range = 0s, 60s ;
		Average_Cloud_Pixel_Distance_Land_Ocean:_FillValue = -9999s ;
		Average_Cloud_Pixel_Distance_Land_Ocean:long_name = "Average Distance (number of pixels) to nearest pixel identified as cloudy from each clear pixel used for Aerosol Retrieval in 10 km retrieval box" ; 
		Average_Cloud_Pixel_Distance_Land_Ocean:units = "Number of Pixels" ;
		Average_Cloud_Pixel_Distance_Land_Ocean:scale_factor = 1. ;
		Average_Cloud_Pixel_Distance_Land_Ocean:add_offset = 0. ;
		Average_Cloud_Pixel_Distance_Land_Ocean:Parameter_Type = "Output" ;
		Average_Cloud_Pixel_Distance_Land_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Average_Cloud_Pixel_Distance_Land_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Average_Cloud_Pixel_Distance_Land_Ocean:_Storage = "chunked" ;
        Average_Cloud_Pixel_Distance_Land_Ocean:_ChunkSizes = 1, 400 ;
        Average_Cloud_Pixel_Distance_Land_Ocean:_DeflateLevel = 5 ;
        Average_Cloud_Pixel_Distance_Land_Ocean:_Shuffle = "true" ;
	short Land_Ocean_Quality_Flag(number_of_lines_8x8, number_of_pixels_8x8) ;
		Land_Ocean_Quality_Flag:valid_range = 0s, 3s ;
		Land_Ocean_Quality_Flag:_FillValue = -9999s ;
		Land_Ocean_Quality_Flag:long_name = "Quality flag for land and ocean aerosol retrievals 0 = Bad  1 = Marginal 2 = Good 3 = Very Good)" ;
		Land_Ocean_Quality_Flag:units = "None" ;
		Land_Ocean_Quality_Flag:scale_factor = 1. ;
		Land_Ocean_Quality_Flag:add_offset = 0. ;
		Land_Ocean_Quality_Flag:Parameter_Type = "Output" ;
		Land_Ocean_Quality_Flag:Geolocation_Pointer = "Internal geolocation arrays" ;
		Land_Ocean_Quality_Flag:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Land_Ocean_Quality_Flag:_Storage = "chunked" ;
        Land_Ocean_Quality_Flag:_ChunkSizes = 1, 400 ;
        Land_Ocean_Quality_Flag:_DeflateLevel = 5 ;
        Land_Ocean_Quality_Flag:_Shuffle = "true" ;
	short Optical_Depth_Land_And_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Optical_Depth_Land_And_Ocean:valid_range = -50s, 5000s ;
		Optical_Depth_Land_And_Ocean:_FillValue = -9999s ;
		Optical_Depth_Land_And_Ocean:long_name = "AOT at 0.55 micron for both ocean (Average) (Quality flag = 1, 2, 3) and land (corrected) (Quality flag = 3)" ;
		Optical_Depth_Land_And_Ocean:units = "None" ;
		Optical_Depth_Land_And_Ocean:scale_factor = 0.001 ;
		Optical_Depth_Land_And_Ocean:add_offset = 0. ;
		Optical_Depth_Land_And_Ocean:Parameter_Type = "Output" ;
		Optical_Depth_Land_And_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Land_And_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Optical_Depth_Land_And_Ocean:_Storage = "chunked" ;
        Optical_Depth_Land_And_Ocean:_ChunkSizes = 1, 400 ;
        Optical_Depth_Land_And_Ocean:_DeflateLevel = 5 ;
        Optical_Depth_Land_And_Ocean:_Shuffle = "true" ;
	short Image_Optical_Depth_Land_And_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Image_Optical_Depth_Land_And_Ocean:valid_range = -50s, 5000s ;
		Image_Optical_Depth_Land_And_Ocean:_FillValue = -9999s ;
		Image_Optical_Depth_Land_And_Ocean:long_name = "AOT at 0.55 micron for both ocean (Average) and land (corrected) with all quality data (Quality flag = 0, 1, 2, 3)" ;
		Image_Optical_Depth_Land_And_Ocean:units = "None" ;
		Image_Optical_Depth_Land_And_Ocean:scale_factor = 0.001 ;
		Image_Optical_Depth_Land_And_Ocean:add_offset = 0. ;
		Image_Optical_Depth_Land_And_Ocean:Parameter_Type = "Output" ;
		Image_Optical_Depth_Land_And_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Image_Optical_Depth_Land_And_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Image_Optical_Depth_Land_And_Ocean:_Storage = "chunked" ;
        Image_Optical_Depth_Land_And_Ocean:_ChunkSizes = 1, 400 ;
        Image_Optical_Depth_Land_And_Ocean:_DeflateLevel = 5 ;
        Image_Optical_Depth_Land_And_Ocean:_Shuffle = "true" ;
	short Aerosol_Type_Land(number_of_lines_8x8, number_of_pixels_8x8) ;
		Aerosol_Type_Land:valid_range = 0s, 4s ;
		Aerosol_Type_Land:_FillValue = -9999s ;
		Aerosol_Type_Land:long_name = "Aerosol Type: 1 = Continental, 2 = Moderate Absorption Fine, 3 = Strong Absorption Fine, 4 = Weak Absorption Fine, 5 = Dust Coarse" ;
		Aerosol_Type_Land:units = "None" ;
		Aerosol_Type_Land:scale_factor = 1. ;
		Aerosol_Type_Land:add_offset = 0. ;
		Aerosol_Type_Land:Parameter_Type = "Output" ;
		Aerosol_Type_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Aerosol_Type_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Aerosol_Type_Land:_Storage = "chunked" ;
        Aerosol_Type_Land:_ChunkSizes = 1, 400 ;
        Aerosol_Type_Land:_DeflateLevel = 5 ;
        Aerosol_Type_Land:_Shuffle = "true" ;
	short Fitting_Error_Land(number_of_lines_8x8, number_of_pixels_8x8) ;
		Fitting_Error_Land:valid_range = 0s, 1000s ;
		Fitting_Error_Land:_FillValue = -9999s ;
		Fitting_Error_Land:long_name = "Spectral Fitting Error for inversion over land" ;
		Fitting_Error_Land:units = "None" ;
		Fitting_Error_Land:scale_factor = 0.001 ;
		Fitting_Error_Land:add_offset = 0. ;
		Fitting_Error_Land:Parameter_Type = "Output" ;
		Fitting_Error_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Fitting_Error_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Fitting_Error_Land:_Storage = "chunked" ;
        Fitting_Error_Land:_ChunkSizes = 1, 400 ;
        Fitting_Error_Land:_DeflateLevel = 5 ;
        Fitting_Error_Land:_Shuffle = "true" ;
	short Surface_Reflectance_Land(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Land_1) ;
		Surface_Reflectance_Land:valid_range = 0s, 1000s ;
		Surface_Reflectance_Land:_FillValue = -9999s ;
		Surface_Reflectance_Land:long_name = "Estimated Surface Reflectance at 0.48, 0.67, 2.25 microns" ;
		Surface_Reflectance_Land:units = "None" ;
		Surface_Reflectance_Land:scale_factor = 0.001 ;
		Surface_Reflectance_Land:add_offset = 0. ;
		Surface_Reflectance_Land:Parameter_Type = "Output" ;
		Surface_Reflectance_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Surface_Reflectance_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude " ;
        Surface_Reflectance_Land:_Storage = "chunked" ;
        Surface_Reflectance_Land:_ChunkSizes = 1, 400, 3 ;
        Surface_Reflectance_Land:_DeflateLevel = 5 ;
        Surface_Reflectance_Land:_Shuffle = "true" ;
	short Corrected_Optical_Depth_Land(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Land_2) ;
		Corrected_Optical_Depth_Land:valid_range = -50s, 5000s ;
		Corrected_Optical_Depth_Land:_FillValue = -9999s ;
		Corrected_Optical_Depth_Land:long_name = "Retrieved AOT at 0.48, 0.55, 0.67, 2.25 microns" ;
		Corrected_Optical_Depth_Land:units = "None" ;
		Corrected_Optical_Depth_Land:scale_factor = 0.001 ;
		Corrected_Optical_Depth_Land:add_offset = 0. ;
		Corrected_Optical_Depth_Land:Parameter_Type = "Output" ;
		Corrected_Optical_Depth_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Corrected_Optical_Depth_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude " ;
        Corrected_Optical_Depth_Land:_Storage = "chunked" ;
        Corrected_Optical_Depth_Land:_ChunkSizes = 1, 400, 4 ;
        Corrected_Optical_Depth_Land:_DeflateLevel = 5 ;
        Corrected_Optical_Depth_Land:_Shuffle = "true" ;
	short Optical_Depth_Ratio_Small_Land(number_of_lines_8x8, number_of_pixels_8x8) ;
		Optical_Depth_Ratio_Small_Land:valid_range = 0s, 1000s ;
		Optical_Depth_Ratio_Small_Land:_FillValue = -9999s ;
		Optical_Depth_Ratio_Small_Land:long_name = "Fraction of AOT contributed by fine dominated model" ;
		Optical_Depth_Ratio_Small_Land:units = "None" ;
		Optical_Depth_Ratio_Small_Land:scale_factor = 0.001 ;
		Optical_Depth_Ratio_Small_Land:add_offset = 0. ;
		Optical_Depth_Ratio_Small_Land:Parameter_Type = "Output" ;
		Optical_Depth_Ratio_Small_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Ratio_Small_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Optical_Depth_Ratio_Small_Land:_Storage = "chunked" ;
        Optical_Depth_Ratio_Small_Land:_ChunkSizes = 1, 400 ;
        Optical_Depth_Ratio_Small_Land:_DeflateLevel = 5 ;
        Optical_Depth_Ratio_Small_Land:_Shuffle = "true" ;
	short Number_Pixels_Used_Land(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Land_1) ;
		Number_Pixels_Used_Land:valid_range = 1s, 400s ;
		Number_Pixels_Used_Land:_FillValue = -9999s ;
		Number_Pixels_Used_Land:long_name = "Number of pixels used for land retrieval at 0.48, 0.67, 2.25 microns" ;
		Number_Pixels_Used_Land:units = "None" ;
		Number_Pixels_Used_Land:scale_factor = 1. ;
		Number_Pixels_Used_Land:add_offset = 0. ;
		Number_Pixels_Used_Land:Parameter_Type = "Output" ;
		Number_Pixels_Used_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Number_Pixels_Used_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Number_Pixels_Used_Land:_Storage = "chunked" ;
        Number_Pixels_Used_Land:_ChunkSizes = 1, 400, 3 ;
        Number_Pixels_Used_Land:_DeflateLevel = 5 ;
        Number_Pixels_Used_Land:_Shuffle = "true" ;
	short Mean_Reflectance_Land(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Land_1) ;
		Mean_Reflectance_Land:valid_range = 0s, 10000s ;
		Mean_Reflectance_Land:_FillValue = -9999s ;
		Mean_Reflectance_Land:long_name = "Mean reflectance of pixels used for land retrieval at 0.48, 0.67, 2.25 microns" ;
		Mean_Reflectance_Land:units = "None" ;
		Mean_Reflectance_Land:scale_factor = 0.0001 ;
		Mean_Reflectance_Land:add_offset = 0. ;
		Mean_Reflectance_Land:Parameter_Type = "Output" ;
		Mean_Reflectance_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mean_Reflectance_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Mean_Reflectance_Land:_Storage = "chunked" ;
        Mean_Reflectance_Land:_ChunkSizes = 1, 400, 3 ;
        Mean_Reflectance_Land:_DeflateLevel = 5 ;
        Mean_Reflectance_Land:_Shuffle = "true" ;
	short STD_Reflectance_Land(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Land_1) ;
		STD_Reflectance_Land:valid_range = 0s, 20000s ;
		STD_Reflectance_Land:_FillValue = -9999s ;
		STD_Reflectance_Land:long_name = "Standard deviation of reflectance of pixels used for land retrieval used for land retrieval at 0.48, 0.67, 2.25 microns" ;
		STD_Reflectance_Land:units = "None" ;
		STD_Reflectance_Land:scale_factor = 0.0001 ;
		STD_Reflectance_Land:add_offset = 0. ;
		STD_Reflectance_Land:Parameter_Type = "Output" ;
		STD_Reflectance_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		STD_Reflectance_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        STD_Reflectance_Land:_Storage = "chunked" ;
        STD_Reflectance_Land:_ChunkSizes = 1, 400, 3 ;
        STD_Reflectance_Land:_DeflateLevel = 5 ;
        STD_Reflectance_Land:_Shuffle = "true" ;
	float Mass_Concentration_Land(number_of_lines_8x8, number_of_pixels_8x8) ;
		Mass_Concentration_Land:valid_range = 0.f, 1000.f ;
		Mass_Concentration_Land:_FillValue = -999.f ;
		Mass_Concentration_Land:long_name = "Estimated Column Mass(per area) using assumed mass extinction efficiency" ;
		Mass_Concentration_Land:units = "1.0e-6g/cm^2" ;
		Mass_Concentration_Land:scale_factor = 1. ;
		Mass_Concentration_Land:add_offset = 0. ;
		Mass_Concentration_Land:Parameter_Type = "Output" ;
		Mass_Concentration_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mass_Concentration_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Mass_Concentration_Land:_Storage = "chunked" ;
        Mass_Concentration_Land:_ChunkSizes = 1, 400 ;
        Mass_Concentration_Land:_DeflateLevel = 5 ;
        Mass_Concentration_Land:_Shuffle = "true" ;
	short Aerosol_Cloud_Fraction_Land(number_of_lines_8x8, number_of_pixels_8x8) ;
		Aerosol_Cloud_Fraction_Land:valid_range = 0s, 1000s ;
		Aerosol_Cloud_Fraction_Land:_FillValue = -9999s ;
		Aerosol_Cloud_Fraction_Land:long_name = "Cloud fraction from Land aerosol cloud mask from retrieved and overcast pixels not including cirrus mask" ;
		Aerosol_Cloud_Fraction_Land:units = "None" ;
		Aerosol_Cloud_Fraction_Land:scale_factor = 0.001 ;
		Aerosol_Cloud_Fraction_Land:add_offset = 0. ;
		Aerosol_Cloud_Fraction_Land:Parameter_Type = "Output" ;
		Aerosol_Cloud_Fraction_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Aerosol_Cloud_Fraction_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Aerosol_Cloud_Fraction_Land:_Storage = "chunked" ;
        Aerosol_Cloud_Fraction_Land:_ChunkSizes = 1, 400 ;
        Aerosol_Cloud_Fraction_Land:_DeflateLevel = 5 ;
        Aerosol_Cloud_Fraction_Land:_Shuffle = "true" ;
	short Effective_Optical_Depth_Average_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		Effective_Optical_Depth_Average_Ocean:valid_range = -50s, 5000s ;
		Effective_Optical_Depth_Average_Ocean:_FillValue = -9999s ;
		Effective_Optical_Depth_Average_Ocean:long_name = "Retrieved AOT for average solution at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Effective_Optical_Depth_Average_Ocean:units = "None" ;
		Effective_Optical_Depth_Average_Ocean:scale_factor = 0.001 ;
		Effective_Optical_Depth_Average_Ocean:add_offset = 0. ;
		Effective_Optical_Depth_Average_Ocean:Parameter_Type = "Output" ;
		Effective_Optical_Depth_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Effective_Optical_Depth_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Effective_Optical_Depth_Average_Ocean:_Storage = "chunked" ;
        Effective_Optical_Depth_Average_Ocean:_ChunkSizes = 1, 400, 7 ;
        Effective_Optical_Depth_Average_Ocean:_DeflateLevel = 5 ;
        Effective_Optical_Depth_Average_Ocean:_Shuffle = "true" ;
	short Optical_Depth_Small_Average_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		Optical_Depth_Small_Average_Ocean:valid_range = -50s, 5000s ;
		Optical_Depth_Small_Average_Ocean:_FillValue = -9999s ;
		Optical_Depth_Small_Average_Ocean:long_name = "Retrieved optical thickness for fine mode (Average solution) for 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Optical_Depth_Small_Average_Ocean:units = "None" ;
		Optical_Depth_Small_Average_Ocean:scale_factor = 0.001 ;
		Optical_Depth_Small_Average_Ocean:add_offset = 0. ;
		Optical_Depth_Small_Average_Ocean:Parameter_Type = "Output" ;
		Optical_Depth_Small_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Small_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Optical_Depth_Small_Average_Ocean:_Storage = "chunked" ;
        Optical_Depth_Small_Average_Ocean:_ChunkSizes = 1, 400, 7 ;
        Optical_Depth_Small_Average_Ocean:_DeflateLevel = 5 ;
        Optical_Depth_Small_Average_Ocean:_Shuffle = "true" ;
	short Optical_Depth_Large_Average_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		Optical_Depth_Large_Average_Ocean:valid_range = -50s, 5000s ;
		Optical_Depth_Large_Average_Ocean:_FillValue = -9999s ;
		Optical_Depth_Large_Average_Ocean:long_name = "Retrieved AOT of large mode for  average  solution at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Optical_Depth_Large_Average_Ocean:units = "None" ;
		Optical_Depth_Large_Average_Ocean:scale_factor = 0.001 ;
		Optical_Depth_Large_Average_Ocean:add_offset = 0. ;
		Optical_Depth_Large_Average_Ocean:Parameter_Type = "Output" ;
		Optical_Depth_Large_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Large_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Optical_Depth_Large_Average_Ocean:_Storage = "chunked" ;
        Optical_Depth_Large_Average_Ocean:_ChunkSizes = 1, 400, 7 ;
        Optical_Depth_Large_Average_Ocean:_DeflateLevel = 5 ;
        Optical_Depth_Large_Average_Ocean:_Shuffle = "true" ;
	float Mass_Concentration_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Mass_Concentration_Ocean:valid_range = 0.f, 1000.f ;
		Mass_Concentration_Ocean:_FillValue = -999.f ;
		Mass_Concentration_Ocean:long_name = "Estimated Column Mass (per area) using assumed mass extinction coefficients" ;
		Mass_Concentration_Ocean:units = "1.0e-6g/cm^2" ;
		Mass_Concentration_Ocean:scale_factor = 1. ;
		Mass_Concentration_Ocean:add_offset = 0. ;
		Mass_Concentration_Ocean:Parameter_Type = "Output" ;
		Mass_Concentration_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mass_Concentration_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Mass_Concentration_Ocean:_Storage = "chunked" ;
        Mass_Concentration_Ocean:_ChunkSizes = 1, 400 ;
        Mass_Concentration_Ocean:_DeflateLevel = 5 ;
        Mass_Concentration_Ocean:_Shuffle = "true" ;
	short Aerosol_Cloud_Fraction_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Aerosol_Cloud_Fraction_Ocean:valid_range = 0s, 1000s ;
		Aerosol_Cloud_Fraction_Ocean:_FillValue = -9999s ;
		Aerosol_Cloud_Fraction_Ocean:long_name = "Cloud fraction from Ocean aerosol cloud mask from retrieved and overcast pixels not including cirrus mask" ;
		Aerosol_Cloud_Fraction_Ocean:units = "None" ;
		Aerosol_Cloud_Fraction_Ocean:scale_factor = 0.001 ;
		Aerosol_Cloud_Fraction_Ocean:add_offset = 0. ;
		Aerosol_Cloud_Fraction_Ocean:Parameter_Type = "Output" ;
		Aerosol_Cloud_Fraction_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Aerosol_Cloud_Fraction_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Aerosol_Cloud_Fraction_Ocean:_Storage = "chunked" ;
        Aerosol_Cloud_Fraction_Ocean:_ChunkSizes = 1, 400 ;
        Aerosol_Cloud_Fraction_Ocean:_DeflateLevel = 5 ;
        Aerosol_Cloud_Fraction_Ocean:_Shuffle = "true" ;
	short Effective_Radius_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Effective_Radius_Ocean:valid_range = 0s, 5000s ;
		Effective_Radius_Ocean:_FillValue = -9999s ;
		Effective_Radius_Ocean:long_name = "Effective_Radius at 0.55 microns" ;
		Effective_Radius_Ocean:units = "micron" ;
		Effective_Radius_Ocean:scale_factor = 0.001 ;
		Effective_Radius_Ocean:add_offset = 0. ;
		Effective_Radius_Ocean:Parameter_Type = "Output" ;
		Effective_Radius_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Effective_Radius_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Effective_Radius_Ocean:_Storage = "chunked" ;
        Effective_Radius_Ocean:_ChunkSizes = 1, 400 ;
        Effective_Radius_Ocean:_DeflateLevel = 5 ;
        Effective_Radius_Ocean:_Shuffle = "true" ;
	float PSML003_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		PSML003_Ocean:valid_range = 0.f, 9.9999998e+10f ;
		PSML003_Ocean:_FillValue = -999.f ;
		PSML003_Ocean:long_name = "Inferred column number concentration (number per area) of particles larger than 0.03 microns" ;
		PSML003_Ocean:units = "Particles/cm^2" ;
		PSML003_Ocean:scale_factor = 1. ;
		PSML003_Ocean:add_offset = 0. ;
		PSML003_Ocean:Parameter_Type = "Output" ;
		PSML003_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		PSML003_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        PSML003_Ocean:_Storage = "chunked" ;
        PSML003_Ocean:_ChunkSizes = 1, 400 ;
        PSML003_Ocean:_DeflateLevel = 5 ;
        PSML003_Ocean:_Shuffle = "true" ;
	short Asymmetry_Factor_Average_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		Asymmetry_Factor_Average_Ocean:valid_range = 0s, 3000s ;
		Asymmetry_Factor_Average_Ocean:_FillValue = -9999s ;
		Asymmetry_Factor_Average_Ocean:long_name = "Inferred Asymmetry_Factor for average solution at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Asymmetry_Factor_Average_Ocean:units = "None" ;
		Asymmetry_Factor_Average_Ocean:scale_factor = 0.001 ;
		Asymmetry_Factor_Average_Ocean:add_offset = 0. ;
		Asymmetry_Factor_Average_Ocean:Parameter_Type = "Output" ;
		Asymmetry_Factor_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Asymmetry_Factor_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Asymmetry_Factor_Average_Ocean:_Storage = "chunked" ;
        Asymmetry_Factor_Average_Ocean:_ChunkSizes = 1, 400, 7 ;
        Asymmetry_Factor_Average_Ocean:_DeflateLevel = 5 ;
        Asymmetry_Factor_Average_Ocean:_Shuffle = "true" ;
	short Backscattering_Ratio_Average_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		Backscattering_Ratio_Average_Ocean:valid_range = 0s, 3000s ;
		Backscattering_Ratio_Average_Ocean:_FillValue = -9999s ;
		Backscattering_Ratio_Average_Ocean:long_name = "Inferred Backscattering Ratio for average solution at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Backscattering_Ratio_Average_Ocean:units = "None" ;
		Backscattering_Ratio_Average_Ocean:scale_factor = 0.001 ;
		Backscattering_Ratio_Average_Ocean:add_offset = 0. ;
		Backscattering_Ratio_Average_Ocean:Parameter_Type = "Output" ;
		Backscattering_Ratio_Average_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Backscattering_Ratio_Average_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Backscattering_Ratio_Average_Ocean:_Storage = "chunked" ;
        Backscattering_Ratio_Average_Ocean:_ChunkSizes = 1, 400, 7 ;
        Backscattering_Ratio_Average_Ocean:_DeflateLevel = 5 ;
        Backscattering_Ratio_Average_Ocean:_Shuffle = "true" ;
	short Angstrom_Exponent_1_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Angstrom_Exponent_1_Ocean:valid_range = -1000s, 5000s ;
		Angstrom_Exponent_1_Ocean:_FillValue = -9999s ;
		Angstrom_Exponent_1_Ocean:long_name = "Calculated Angstrom Exponent for 0.55 vs 0.86 micron for Average Solution" ;
		Angstrom_Exponent_1_Ocean:units = "None" ;
		Angstrom_Exponent_1_Ocean:scale_factor = 0.001 ;
		Angstrom_Exponent_1_Ocean:add_offset = 0. ;
		Angstrom_Exponent_1_Ocean:Parameter_Type = "Output" ;
		Angstrom_Exponent_1_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Angstrom_Exponent_1_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Angstrom_Exponent_1_Ocean:_Storage = "chunked" ;
        Angstrom_Exponent_1_Ocean:_ChunkSizes = 1, 400 ;
        Angstrom_Exponent_1_Ocean:_DeflateLevel = 5 ;
        Angstrom_Exponent_1_Ocean:_Shuffle = "true" ;
	short Angstrom_Exponent_2_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Angstrom_Exponent_2_Ocean:valid_range = -1000s, 5000s ;
		Angstrom_Exponent_2_Ocean:_FillValue = -9999s ;
		Angstrom_Exponent_2_Ocean:long_name = "Calculated Angstrom Exponent for 0.86 vs 2.13 micron for Average Solution" ;
		Angstrom_Exponent_2_Ocean:units = "None" ;
		Angstrom_Exponent_2_Ocean:scale_factor = 0.001 ;
		Angstrom_Exponent_2_Ocean:add_offset = 0. ;
		Angstrom_Exponent_2_Ocean:Parameter_Type = "Output" ;
		Angstrom_Exponent_2_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Angstrom_Exponent_2_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Angstrom_Exponent_2_Ocean:_Storage = "chunked" ;
        Angstrom_Exponent_2_Ocean:_ChunkSizes = 1, 400 ;
        Angstrom_Exponent_2_Ocean:_DeflateLevel = 5 ;
        Angstrom_Exponent_2_Ocean:_Shuffle = "true" ;
	short Least_Squares_Error_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Least_Squares_Error_Ocean:valid_range = 0s, 1000s ;
		Least_Squares_Error_Ocean:_FillValue = -9999s ;
		Least_Squares_Error_Ocean:long_name = "Residual of least squares fitting for inversion over ocean" ;
		Least_Squares_Error_Ocean:units = "None" ;
		Least_Squares_Error_Ocean:scale_factor = 0.001 ;
		Least_Squares_Error_Ocean:add_offset = 0. ;
		Least_Squares_Error_Ocean:Parameter_Type = "Output" ;
		Least_Squares_Error_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Least_Squares_Error_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Least_Squares_Error_Ocean:_Storage = "chunked" ;
        Least_Squares_Error_Ocean:_ChunkSizes = 1, 400 ;
        Least_Squares_Error_Ocean:_DeflateLevel = 5 ;
        Least_Squares_Error_Ocean:_Shuffle = "true" ;
	short Optical_Depth_Ratio_Small_Ocean_0p55micron(number_of_lines_8x8, number_of_pixels_8x8) ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:valid_range = 0s, 1000s ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:_FillValue = -9999s ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:long_name = "Fraction of AOT (at 0.55 micron) contributed by fine mode for average solution" ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:units = "None" ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:scale_factor = 0.001 ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:add_offset = 0. ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:Parameter_Type = "Output" ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_Ratio_Small_Ocean_0p55micron:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Optical_Depth_Ratio_Small_Ocean_0p55micron:_Storage = "chunked" ;
        Optical_Depth_Ratio_Small_Ocean_0p55micron:_ChunkSizes = 1, 400 ;
        Optical_Depth_Ratio_Small_Ocean_0p55micron:_DeflateLevel = 5 ;
        Optical_Depth_Ratio_Small_Ocean_0p55micron:_Shuffle = "true" ;
	short Optical_Depth_By_Models_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Solution_Index) ;
		Optical_Depth_By_Models_Ocean:valid_range = -50s, 5000s ;
		Optical_Depth_By_Models_Ocean:_FillValue = -9999s ;
		Optical_Depth_By_Models_Ocean:long_name = "Retrieved AOT (at 0.55 micron) partioned by mode index (for Best solution)" ;
		Optical_Depth_By_Models_Ocean:units = "None" ;
		Optical_Depth_By_Models_Ocean:scale_factor = 0.001 ;
		Optical_Depth_By_Models_Ocean:add_offset = 0. ;
		Optical_Depth_By_Models_Ocean:Parameter_Type = "Output" ;
		Optical_Depth_By_Models_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Optical_Depth_By_Models_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Optical_Depth_By_Models_Ocean:_Storage = "chunked" ;
        Optical_Depth_By_Models_Ocean:_ChunkSizes = 1, 400, 9 ;
        Optical_Depth_By_Models_Ocean:_DeflateLevel = 5 ;
        Optical_Depth_By_Models_Ocean:_Shuffle = "true" ;
	short Number_Pixels_Used_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		Number_Pixels_Used_Ocean:valid_range = 1s, 400s ;
		Number_Pixels_Used_Ocean:_FillValue = -9999s ;
		Number_Pixels_Used_Ocean:long_name = "Number of pixels used for ocean retrieval at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Number_Pixels_Used_Ocean:units = "None" ;
		Number_Pixels_Used_Ocean:scale_factor = 1. ;
		Number_Pixels_Used_Ocean:add_offset = 0. ;
		Number_Pixels_Used_Ocean:Parameter_Type = "Output" ;
		Number_Pixels_Used_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Number_Pixels_Used_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Number_Pixels_Used_Ocean:_Storage = "chunked" ;
        Number_Pixels_Used_Ocean:_ChunkSizes = 1, 400, 7 ;
        Number_Pixels_Used_Ocean:_DeflateLevel = 5 ;
        Number_Pixels_Used_Ocean:_Shuffle = "true" ;
	short Mean_Reflectance_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		Mean_Reflectance_Ocean:valid_range = 0s, 10000s ;
		Mean_Reflectance_Ocean:_FillValue = -9999s ;
		Mean_Reflectance_Ocean:long_name = "Mean reflectance of pixels used for ocean retrieval at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		Mean_Reflectance_Ocean:units = "None" ;
		Mean_Reflectance_Ocean:scale_factor = 0.0001 ;
		Mean_Reflectance_Ocean:add_offset = 0. ;
		Mean_Reflectance_Ocean:Parameter_Type = "Output" ;
		Mean_Reflectance_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Mean_Reflectance_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Mean_Reflectance_Ocean:_Storage = "chunked" ;
        Mean_Reflectance_Ocean:_ChunkSizes = 1, 400, 7 ;
        Mean_Reflectance_Ocean:_DeflateLevel = 5 ;
        Mean_Reflectance_Ocean:_Shuffle = "true" ;
	short STD_Reflectance_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Wavelength_Used_Ocean) ;
		STD_Reflectance_Ocean:valid_range = 0s, 20000s ;
		STD_Reflectance_Ocean:_FillValue = -9999s ;
		STD_Reflectance_Ocean:long_name = "Standard deviation of reflectance of pixels used for ocean retrieval at 0.48, 0.55, 0.67, 0.86, 1.24, 1.60, 2.25 microns" ;
		STD_Reflectance_Ocean:units = "None" ;
		STD_Reflectance_Ocean:scale_factor = 0.0001 ;
		STD_Reflectance_Ocean:add_offset = 0. ;
		STD_Reflectance_Ocean:Parameter_Type = "Output" ;
		STD_Reflectance_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		STD_Reflectance_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        STD_Reflectance_Ocean:_Storage = "chunked" ;
        STD_Reflectance_Ocean:_ChunkSizes = 1, 400, 7 ;
        STD_Reflectance_Ocean:_DeflateLevel = 5 ;
        STD_Reflectance_Ocean:_Shuffle = "true" ;
	short Wind_Speed_Ncep_Ocean(number_of_lines_8x8, number_of_pixels_8x8) ;
		Wind_Speed_Ncep_Ocean:valid_range = 0s, 8000s ;
		Wind_Speed_Ncep_Ocean:_FillValue = -9999s ;
		Wind_Speed_Ncep_Ocean:long_name = "Wind Speed based on NCEP reanalysis for Ocean" ;
		Wind_Speed_Ncep_Ocean:units = "Meters/sec" ;
		Wind_Speed_Ncep_Ocean:scale_factor = 0.01 ;
		Wind_Speed_Ncep_Ocean:add_offset = 0. ;
		Wind_Speed_Ncep_Ocean:Parameter_Type = "Output" ;
		Wind_Speed_Ncep_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Wind_Speed_Ncep_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Wind_Speed_Ncep_Ocean:_Storage = "chunked" ;
        Wind_Speed_Ncep_Ocean:_ChunkSizes = 1, 400 ;
        Wind_Speed_Ncep_Ocean:_DeflateLevel = 5 ;
        Wind_Speed_Ncep_Ocean:_Shuffle = "true" ;
	short Topographic_Altitude_Land(number_of_lines_8x8, number_of_pixels_8x8) ;
		Topographic_Altitude_Land:valid_range = 0s, 1000s ;
		Topographic_Altitude_Land:_FillValue = -9999s ;
		Topographic_Altitude_Land:long_name = "Averaged topographic altitude (in km) for Land" ;
		Topographic_Altitude_Land:units = "KM" ;
		Topographic_Altitude_Land:scale_factor = 0.01 ;
		Topographic_Altitude_Land:add_offset = 0. ;
		Topographic_Altitude_Land:Parameter_Type = "Output" ;
		Topographic_Altitude_Land:Geolocation_Pointer = "Internal geolocation arrays" ;
		Topographic_Altitude_Land:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Topographic_Altitude_Land:_Storage = "chunked" ;
        Topographic_Altitude_Land:_ChunkSizes = 1, 400 ;
        Topographic_Altitude_Land:_DeflateLevel = 5 ;
        Topographic_Altitude_Land:_Shuffle = "true" ;
	short Error_Flag_Land_And_Ocean(number_of_lines_8x8, number_of_pixels_8x8, Quality_Flag_Num) ;
		Error_Flag_Land_And_Ocean:valid_range = 1s, 26s ;
        Error_Flag_Land_And_Ocean:_FillValue = -9999s ;
        Error_Flag_Land_And_Ocean:long_name = "Error code 1-26. Layer 1 ocean, Layer 2 land. Ask for Documentation" ;
        Error_Flag_Land_And_Ocean:units = "None" ;
        Error_Flag_Land_And_Ocean:scale_factor = 1.0 ;
        Error_Flag_Land_And_Ocean:add_offset = 0. ;
        Error_Flag_Land_And_Ocean:Parameter_Type = "Output" ;
        Error_Flag_Land_And_Ocean:Geolocation_Pointer = "Internal geolocation arrays" ;
		Error_Flag_Land_And_Ocean:coordinates = "/geolocation_data/longitude /geolocation_data/latitude" ;
        Error_Flag_Land_And_Ocean:_Storage = "chunked" ;
        Error_Flag_Land_And_Ocean:_ChunkSizes = 1, 400, 2 ;
        Error_Flag_Land_And_Ocean:_DeflateLevel = 5 ;
        Error_Flag_Land_And_Ocean:_Shuffle = "true" ;
    data:
    } // group geophysical_data
}
